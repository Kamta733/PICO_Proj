magic
tech sky130A
magscale 1 2
timestamp 1661836425
<< nwell >>
rect 3530 -2341 9992 2305
<< pwell >>
rect -116 2210 -74 2211
rect -1607 2117 1607 2210
rect -1608 2021 1607 2117
rect -1607 -2210 1607 2021
<< nmos >>
rect -1407 -2000 -1377 2000
rect -1311 -2000 -1281 2000
rect -1215 -2000 -1185 2000
rect -1119 -2000 -1089 2000
rect -1023 -2000 -993 2000
rect -927 -2000 -897 2000
rect -831 -2000 -801 2000
rect -735 -2000 -705 2000
rect -639 -2000 -609 2000
rect -543 -2000 -513 2000
rect -447 -2000 -417 2000
rect -351 -2000 -321 2000
rect -255 -2000 -225 2000
rect -159 -2000 -129 2000
rect -63 -2000 -33 2000
rect 33 -2000 63 2000
rect 129 -2000 159 2000
rect 225 -2000 255 2000
rect 321 -2000 351 2000
rect 417 -2000 447 2000
rect 513 -2000 543 2000
rect 609 -2000 639 2000
rect 705 -2000 735 2000
rect 801 -2000 831 2000
rect 897 -2000 927 2000
rect 993 -2000 1023 2000
rect 1089 -2000 1119 2000
rect 1185 -2000 1215 2000
rect 1281 -2000 1311 2000
rect 1377 -2000 1407 2000
<< pmos >>
rect 3865 -2050 3895 1950
rect 3961 -2050 3991 1950
rect 4057 -2050 4087 1950
rect 4153 -2050 4183 1950
rect 4249 -2050 4279 1950
rect 4345 -2050 4375 1950
rect 4441 -2050 4471 1950
rect 4537 -2050 4567 1950
rect 4633 -2050 4663 1950
rect 4729 -2050 4759 1950
rect 4825 -2050 4855 1950
rect 4921 -2050 4951 1950
rect 5017 -2050 5047 1950
rect 5113 -2050 5143 1950
rect 5209 -2050 5239 1950
rect 5305 -2050 5335 1950
rect 5401 -2050 5431 1950
rect 5497 -2050 5527 1950
rect 5593 -2050 5623 1950
rect 5689 -2050 5719 1950
rect 5785 -2050 5815 1950
rect 5881 -2050 5911 1950
rect 5977 -2050 6007 1950
rect 6073 -2050 6103 1950
rect 6169 -2050 6199 1950
rect 6265 -2050 6295 1950
rect 6361 -2050 6391 1950
rect 6457 -2050 6487 1950
rect 6553 -2050 6583 1950
rect 6649 -2050 6679 1950
rect 6745 -2050 6775 1950
rect 6841 -2050 6871 1950
rect 6937 -2050 6967 1950
rect 7033 -2050 7063 1950
rect 7129 -2050 7159 1950
rect 7225 -2050 7255 1950
rect 7321 -2050 7351 1950
rect 7417 -2050 7447 1950
rect 7513 -2050 7543 1950
rect 7609 -2050 7639 1950
rect 7705 -2050 7735 1950
rect 7801 -2050 7831 1950
rect 7897 -2050 7927 1950
rect 7993 -2050 8023 1950
rect 8089 -2050 8119 1950
rect 8185 -2050 8215 1950
rect 8281 -2050 8311 1950
rect 8377 -2050 8407 1950
rect 8473 -2050 8503 1950
rect 8569 -2050 8599 1950
rect 8665 -2050 8695 1950
rect 8761 -2050 8791 1950
rect 8857 -2050 8887 1950
rect 8953 -2050 8983 1950
rect 9049 -2050 9079 1950
rect 9145 -2050 9175 1950
rect 9241 -2050 9271 1950
rect 9337 -2050 9367 1950
rect 9433 -2050 9463 1950
rect 9529 -2050 9559 1950
<< ndiff >>
rect -1469 1988 -1407 2000
rect -1469 -1988 -1457 1988
rect -1423 -1988 -1407 1988
rect -1469 -2000 -1407 -1988
rect -1377 1988 -1311 2000
rect -1377 -1988 -1361 1988
rect -1327 -1988 -1311 1988
rect -1377 -2000 -1311 -1988
rect -1281 1988 -1215 2000
rect -1281 -1988 -1265 1988
rect -1231 -1988 -1215 1988
rect -1281 -2000 -1215 -1988
rect -1185 1988 -1119 2000
rect -1185 -1988 -1169 1988
rect -1135 -1988 -1119 1988
rect -1185 -2000 -1119 -1988
rect -1089 1988 -1023 2000
rect -1089 -1988 -1073 1988
rect -1039 -1988 -1023 1988
rect -1089 -2000 -1023 -1988
rect -993 1988 -927 2000
rect -993 -1988 -977 1988
rect -943 -1988 -927 1988
rect -993 -2000 -927 -1988
rect -897 1988 -831 2000
rect -897 -1988 -881 1988
rect -847 -1988 -831 1988
rect -897 -2000 -831 -1988
rect -801 1988 -735 2000
rect -801 -1988 -785 1988
rect -751 -1988 -735 1988
rect -801 -2000 -735 -1988
rect -705 1988 -639 2000
rect -705 -1988 -689 1988
rect -655 -1988 -639 1988
rect -705 -2000 -639 -1988
rect -609 1988 -543 2000
rect -609 -1988 -593 1988
rect -559 -1988 -543 1988
rect -609 -2000 -543 -1988
rect -513 1988 -447 2000
rect -513 -1988 -497 1988
rect -463 -1988 -447 1988
rect -513 -2000 -447 -1988
rect -417 1988 -351 2000
rect -417 -1988 -401 1988
rect -367 -1988 -351 1988
rect -417 -2000 -351 -1988
rect -321 1988 -255 2000
rect -321 -1988 -305 1988
rect -271 -1988 -255 1988
rect -321 -2000 -255 -1988
rect -225 1988 -159 2000
rect -225 -1988 -209 1988
rect -175 -1988 -159 1988
rect -225 -2000 -159 -1988
rect -129 1988 -63 2000
rect -129 -1988 -113 1988
rect -79 -1988 -63 1988
rect -129 -2000 -63 -1988
rect -33 1988 33 2000
rect -33 -1988 -17 1988
rect 17 -1988 33 1988
rect -33 -2000 33 -1988
rect 63 1988 129 2000
rect 63 -1988 79 1988
rect 113 -1988 129 1988
rect 63 -2000 129 -1988
rect 159 1988 225 2000
rect 159 -1988 175 1988
rect 209 -1988 225 1988
rect 159 -2000 225 -1988
rect 255 1988 321 2000
rect 255 -1988 271 1988
rect 305 -1988 321 1988
rect 255 -2000 321 -1988
rect 351 1988 417 2000
rect 351 -1988 367 1988
rect 401 -1988 417 1988
rect 351 -2000 417 -1988
rect 447 1988 513 2000
rect 447 -1988 463 1988
rect 497 -1988 513 1988
rect 447 -2000 513 -1988
rect 543 1988 609 2000
rect 543 -1988 559 1988
rect 593 -1988 609 1988
rect 543 -2000 609 -1988
rect 639 1988 705 2000
rect 639 -1988 655 1988
rect 689 -1988 705 1988
rect 639 -2000 705 -1988
rect 735 1988 801 2000
rect 735 -1988 751 1988
rect 785 -1988 801 1988
rect 735 -2000 801 -1988
rect 831 1988 897 2000
rect 831 -1988 847 1988
rect 881 -1988 897 1988
rect 831 -2000 897 -1988
rect 927 1988 993 2000
rect 927 -1988 943 1988
rect 977 -1988 993 1988
rect 927 -2000 993 -1988
rect 1023 1988 1089 2000
rect 1023 -1988 1039 1988
rect 1073 -1988 1089 1988
rect 1023 -2000 1089 -1988
rect 1119 1988 1185 2000
rect 1119 -1988 1135 1988
rect 1169 -1988 1185 1988
rect 1119 -2000 1185 -1988
rect 1215 1988 1281 2000
rect 1215 -1988 1231 1988
rect 1265 -1988 1281 1988
rect 1215 -2000 1281 -1988
rect 1311 1988 1377 2000
rect 1311 -1988 1327 1988
rect 1361 -1988 1377 1988
rect 1311 -2000 1377 -1988
rect 1407 1988 1469 2000
rect 1407 -1988 1423 1988
rect 1457 -1988 1469 1988
rect 1407 -2000 1469 -1988
<< pdiff >>
rect 3803 1938 3865 1950
rect 3803 -2038 3815 1938
rect 3849 -2038 3865 1938
rect 3803 -2050 3865 -2038
rect 3895 1938 3961 1950
rect 3895 -2038 3911 1938
rect 3945 -2038 3961 1938
rect 3895 -2050 3961 -2038
rect 3991 1938 4057 1950
rect 3991 -2038 4007 1938
rect 4041 -2038 4057 1938
rect 3991 -2050 4057 -2038
rect 4087 1938 4153 1950
rect 4087 -2038 4103 1938
rect 4137 -2038 4153 1938
rect 4087 -2050 4153 -2038
rect 4183 1938 4249 1950
rect 4183 -2038 4199 1938
rect 4233 -2038 4249 1938
rect 4183 -2050 4249 -2038
rect 4279 1938 4345 1950
rect 4279 -2038 4295 1938
rect 4329 -2038 4345 1938
rect 4279 -2050 4345 -2038
rect 4375 1938 4441 1950
rect 4375 -2038 4391 1938
rect 4425 -2038 4441 1938
rect 4375 -2050 4441 -2038
rect 4471 1938 4537 1950
rect 4471 -2038 4487 1938
rect 4521 -2038 4537 1938
rect 4471 -2050 4537 -2038
rect 4567 1938 4633 1950
rect 4567 -2038 4583 1938
rect 4617 -2038 4633 1938
rect 4567 -2050 4633 -2038
rect 4663 1938 4729 1950
rect 4663 -2038 4679 1938
rect 4713 -2038 4729 1938
rect 4663 -2050 4729 -2038
rect 4759 1938 4825 1950
rect 4759 -2038 4775 1938
rect 4809 -2038 4825 1938
rect 4759 -2050 4825 -2038
rect 4855 1938 4921 1950
rect 4855 -2038 4871 1938
rect 4905 -2038 4921 1938
rect 4855 -2050 4921 -2038
rect 4951 1938 5017 1950
rect 4951 -2038 4967 1938
rect 5001 -2038 5017 1938
rect 4951 -2050 5017 -2038
rect 5047 1938 5113 1950
rect 5047 -2038 5063 1938
rect 5097 -2038 5113 1938
rect 5047 -2050 5113 -2038
rect 5143 1938 5209 1950
rect 5143 -2038 5159 1938
rect 5193 -2038 5209 1938
rect 5143 -2050 5209 -2038
rect 5239 1938 5305 1950
rect 5239 -2038 5255 1938
rect 5289 -2038 5305 1938
rect 5239 -2050 5305 -2038
rect 5335 1938 5401 1950
rect 5335 -2038 5351 1938
rect 5385 -2038 5401 1938
rect 5335 -2050 5401 -2038
rect 5431 1938 5497 1950
rect 5431 -2038 5447 1938
rect 5481 -2038 5497 1938
rect 5431 -2050 5497 -2038
rect 5527 1938 5593 1950
rect 5527 -2038 5543 1938
rect 5577 -2038 5593 1938
rect 5527 -2050 5593 -2038
rect 5623 1938 5689 1950
rect 5623 -2038 5639 1938
rect 5673 -2038 5689 1938
rect 5623 -2050 5689 -2038
rect 5719 1938 5785 1950
rect 5719 -2038 5735 1938
rect 5769 -2038 5785 1938
rect 5719 -2050 5785 -2038
rect 5815 1938 5881 1950
rect 5815 -2038 5831 1938
rect 5865 -2038 5881 1938
rect 5815 -2050 5881 -2038
rect 5911 1938 5977 1950
rect 5911 -2038 5927 1938
rect 5961 -2038 5977 1938
rect 5911 -2050 5977 -2038
rect 6007 1938 6073 1950
rect 6007 -2038 6023 1938
rect 6057 -2038 6073 1938
rect 6007 -2050 6073 -2038
rect 6103 1938 6169 1950
rect 6103 -2038 6119 1938
rect 6153 -2038 6169 1938
rect 6103 -2050 6169 -2038
rect 6199 1938 6265 1950
rect 6199 -2038 6215 1938
rect 6249 -2038 6265 1938
rect 6199 -2050 6265 -2038
rect 6295 1938 6361 1950
rect 6295 -2038 6311 1938
rect 6345 -2038 6361 1938
rect 6295 -2050 6361 -2038
rect 6391 1938 6457 1950
rect 6391 -2038 6407 1938
rect 6441 -2038 6457 1938
rect 6391 -2050 6457 -2038
rect 6487 1938 6553 1950
rect 6487 -2038 6503 1938
rect 6537 -2038 6553 1938
rect 6487 -2050 6553 -2038
rect 6583 1938 6649 1950
rect 6583 -2038 6599 1938
rect 6633 -2038 6649 1938
rect 6583 -2050 6649 -2038
rect 6679 1938 6745 1950
rect 6679 -2038 6695 1938
rect 6729 -2038 6745 1938
rect 6679 -2050 6745 -2038
rect 6775 1938 6841 1950
rect 6775 -2038 6791 1938
rect 6825 -2038 6841 1938
rect 6775 -2050 6841 -2038
rect 6871 1938 6937 1950
rect 6871 -2038 6887 1938
rect 6921 -2038 6937 1938
rect 6871 -2050 6937 -2038
rect 6967 1938 7033 1950
rect 6967 -2038 6983 1938
rect 7017 -2038 7033 1938
rect 6967 -2050 7033 -2038
rect 7063 1938 7129 1950
rect 7063 -2038 7079 1938
rect 7113 -2038 7129 1938
rect 7063 -2050 7129 -2038
rect 7159 1938 7225 1950
rect 7159 -2038 7175 1938
rect 7209 -2038 7225 1938
rect 7159 -2050 7225 -2038
rect 7255 1938 7321 1950
rect 7255 -2038 7271 1938
rect 7305 -2038 7321 1938
rect 7255 -2050 7321 -2038
rect 7351 1938 7417 1950
rect 7351 -2038 7367 1938
rect 7401 -2038 7417 1938
rect 7351 -2050 7417 -2038
rect 7447 1938 7513 1950
rect 7447 -2038 7463 1938
rect 7497 -2038 7513 1938
rect 7447 -2050 7513 -2038
rect 7543 1938 7609 1950
rect 7543 -2038 7559 1938
rect 7593 -2038 7609 1938
rect 7543 -2050 7609 -2038
rect 7639 1938 7705 1950
rect 7639 -2038 7655 1938
rect 7689 -2038 7705 1938
rect 7639 -2050 7705 -2038
rect 7735 1938 7801 1950
rect 7735 -2038 7751 1938
rect 7785 -2038 7801 1938
rect 7735 -2050 7801 -2038
rect 7831 1938 7897 1950
rect 7831 -2038 7847 1938
rect 7881 -2038 7897 1938
rect 7831 -2050 7897 -2038
rect 7927 1938 7993 1950
rect 7927 -2038 7943 1938
rect 7977 -2038 7993 1938
rect 7927 -2050 7993 -2038
rect 8023 1938 8089 1950
rect 8023 -2038 8039 1938
rect 8073 -2038 8089 1938
rect 8023 -2050 8089 -2038
rect 8119 1938 8185 1950
rect 8119 -2038 8135 1938
rect 8169 -2038 8185 1938
rect 8119 -2050 8185 -2038
rect 8215 1938 8281 1950
rect 8215 -2038 8231 1938
rect 8265 -2038 8281 1938
rect 8215 -2050 8281 -2038
rect 8311 1938 8377 1950
rect 8311 -2038 8327 1938
rect 8361 -2038 8377 1938
rect 8311 -2050 8377 -2038
rect 8407 1938 8473 1950
rect 8407 -2038 8423 1938
rect 8457 -2038 8473 1938
rect 8407 -2050 8473 -2038
rect 8503 1938 8569 1950
rect 8503 -2038 8519 1938
rect 8553 -2038 8569 1938
rect 8503 -2050 8569 -2038
rect 8599 1938 8665 1950
rect 8599 -2038 8615 1938
rect 8649 -2038 8665 1938
rect 8599 -2050 8665 -2038
rect 8695 1938 8761 1950
rect 8695 -2038 8711 1938
rect 8745 -2038 8761 1938
rect 8695 -2050 8761 -2038
rect 8791 1938 8857 1950
rect 8791 -2038 8807 1938
rect 8841 -2038 8857 1938
rect 8791 -2050 8857 -2038
rect 8887 1938 8953 1950
rect 8887 -2038 8903 1938
rect 8937 -2038 8953 1938
rect 8887 -2050 8953 -2038
rect 8983 1938 9049 1950
rect 8983 -2038 8999 1938
rect 9033 -2038 9049 1938
rect 8983 -2050 9049 -2038
rect 9079 1938 9145 1950
rect 9079 -2038 9095 1938
rect 9129 -2038 9145 1938
rect 9079 -2050 9145 -2038
rect 9175 1938 9241 1950
rect 9175 -2038 9191 1938
rect 9225 -2038 9241 1938
rect 9175 -2050 9241 -2038
rect 9271 1938 9337 1950
rect 9271 -2038 9287 1938
rect 9321 -2038 9337 1938
rect 9271 -2050 9337 -2038
rect 9367 1938 9433 1950
rect 9367 -2038 9383 1938
rect 9417 -2038 9433 1938
rect 9367 -2050 9433 -2038
rect 9463 1938 9529 1950
rect 9463 -2038 9479 1938
rect 9513 -2038 9529 1938
rect 9463 -2050 9529 -2038
rect 9559 1938 9621 1950
rect 9559 -2038 9575 1938
rect 9609 -2038 9621 1938
rect 9559 -2050 9621 -2038
<< ndiffc >>
rect -1457 -1988 -1423 1988
rect -1361 -1988 -1327 1988
rect -1265 -1988 -1231 1988
rect -1169 -1988 -1135 1988
rect -1073 -1988 -1039 1988
rect -977 -1988 -943 1988
rect -881 -1988 -847 1988
rect -785 -1988 -751 1988
rect -689 -1988 -655 1988
rect -593 -1988 -559 1988
rect -497 -1988 -463 1988
rect -401 -1988 -367 1988
rect -305 -1988 -271 1988
rect -209 -1988 -175 1988
rect -113 -1988 -79 1988
rect -17 -1988 17 1988
rect 79 -1988 113 1988
rect 175 -1988 209 1988
rect 271 -1988 305 1988
rect 367 -1988 401 1988
rect 463 -1988 497 1988
rect 559 -1988 593 1988
rect 655 -1988 689 1988
rect 751 -1988 785 1988
rect 847 -1988 881 1988
rect 943 -1988 977 1988
rect 1039 -1988 1073 1988
rect 1135 -1988 1169 1988
rect 1231 -1988 1265 1988
rect 1327 -1988 1361 1988
rect 1423 -1988 1457 1988
<< pdiffc >>
rect 3815 -2038 3849 1938
rect 3911 -2038 3945 1938
rect 4007 -2038 4041 1938
rect 4103 -2038 4137 1938
rect 4199 -2038 4233 1938
rect 4295 -2038 4329 1938
rect 4391 -2038 4425 1938
rect 4487 -2038 4521 1938
rect 4583 -2038 4617 1938
rect 4679 -2038 4713 1938
rect 4775 -2038 4809 1938
rect 4871 -2038 4905 1938
rect 4967 -2038 5001 1938
rect 5063 -2038 5097 1938
rect 5159 -2038 5193 1938
rect 5255 -2038 5289 1938
rect 5351 -2038 5385 1938
rect 5447 -2038 5481 1938
rect 5543 -2038 5577 1938
rect 5639 -2038 5673 1938
rect 5735 -2038 5769 1938
rect 5831 -2038 5865 1938
rect 5927 -2038 5961 1938
rect 6023 -2038 6057 1938
rect 6119 -2038 6153 1938
rect 6215 -2038 6249 1938
rect 6311 -2038 6345 1938
rect 6407 -2038 6441 1938
rect 6503 -2038 6537 1938
rect 6599 -2038 6633 1938
rect 6695 -2038 6729 1938
rect 6791 -2038 6825 1938
rect 6887 -2038 6921 1938
rect 6983 -2038 7017 1938
rect 7079 -2038 7113 1938
rect 7175 -2038 7209 1938
rect 7271 -2038 7305 1938
rect 7367 -2038 7401 1938
rect 7463 -2038 7497 1938
rect 7559 -2038 7593 1938
rect 7655 -2038 7689 1938
rect 7751 -2038 7785 1938
rect 7847 -2038 7881 1938
rect 7943 -2038 7977 1938
rect 8039 -2038 8073 1938
rect 8135 -2038 8169 1938
rect 8231 -2038 8265 1938
rect 8327 -2038 8361 1938
rect 8423 -2038 8457 1938
rect 8519 -2038 8553 1938
rect 8615 -2038 8649 1938
rect 8711 -2038 8745 1938
rect 8807 -2038 8841 1938
rect 8903 -2038 8937 1938
rect 8999 -2038 9033 1938
rect 9095 -2038 9129 1938
rect 9191 -2038 9225 1938
rect 9287 -2038 9321 1938
rect 9383 -2038 9417 1938
rect 9479 -2038 9513 1938
rect 9575 -2038 9609 1938
<< psubdiff >>
rect -1537 -2174 -1473 -2140
rect 1477 -2174 1537 -2140
<< nsubdiff >>
rect 3735 -2224 3799 -2190
rect 9629 -2224 9689 -2190
<< psubdiffcont >>
rect -1473 -2174 1477 -2140
<< nsubdiffcont >>
rect 3799 -2224 9629 -2190
<< poly >>
rect -1584 2071 -1494 2087
rect -1584 2003 -1572 2071
rect -1510 2051 -1494 2071
rect -1510 2021 1462 2051
rect -1510 2003 -1494 2021
rect -1584 1987 -1494 2003
rect -1407 2000 -1377 2021
rect -1311 2000 -1281 2021
rect -1215 2000 -1185 2021
rect -1119 2000 -1089 2021
rect -1023 2000 -993 2021
rect -927 2000 -897 2021
rect -831 2000 -801 2021
rect -735 2000 -705 2021
rect -639 2000 -609 2021
rect -543 2000 -513 2021
rect -447 2000 -417 2021
rect -351 2000 -321 2021
rect -255 2000 -225 2021
rect -159 2000 -129 2021
rect -63 2000 -33 2021
rect 33 2000 63 2021
rect 129 2000 159 2021
rect 225 2000 255 2021
rect 321 2000 351 2021
rect 417 2000 447 2021
rect 513 2000 543 2021
rect 609 2000 639 2021
rect 705 2000 735 2021
rect 801 2000 831 2021
rect 897 2000 927 2021
rect 993 2000 1023 2021
rect 1089 2000 1119 2021
rect 1185 2000 1215 2021
rect 1270 2019 1311 2021
rect 1281 2000 1311 2019
rect 1377 2000 1407 2021
rect 3684 2017 3778 2037
rect 3684 1959 3696 2017
rect 3756 2001 3778 2017
rect 3756 1971 9614 2001
rect 3756 1959 3778 1971
rect 3684 1937 3778 1959
rect 3865 1950 3895 1971
rect 3961 1950 3991 1971
rect 4057 1950 4087 1971
rect 4153 1950 4183 1971
rect 4249 1950 4279 1971
rect 4345 1950 4375 1971
rect 4441 1950 4471 1971
rect 4537 1950 4567 1971
rect 4633 1950 4663 1971
rect 4729 1950 4759 1971
rect 4825 1950 4855 1971
rect 4921 1950 4951 1971
rect 5017 1950 5047 1971
rect 5113 1950 5143 1971
rect 5209 1950 5239 1971
rect 5305 1950 5335 1971
rect 5401 1950 5431 1971
rect 5497 1950 5527 1971
rect 5593 1950 5623 1971
rect 5689 1950 5719 1971
rect 5785 1950 5815 1971
rect 5881 1950 5911 1971
rect 5977 1950 6007 1971
rect 6073 1950 6103 1971
rect 6169 1950 6199 1971
rect 6265 1950 6295 1971
rect 6361 1950 6391 1971
rect 6457 1950 6487 1971
rect 6542 1969 6583 1971
rect 6553 1950 6583 1969
rect 6649 1950 6679 1971
rect 6745 1950 6775 1971
rect 6841 1950 6871 1971
rect 6937 1950 6967 1971
rect 7033 1950 7063 1971
rect 7129 1950 7159 1971
rect 7225 1950 7255 1971
rect 7321 1950 7351 1971
rect 7417 1950 7447 1971
rect 7513 1950 7543 1971
rect 7609 1950 7639 1971
rect 7705 1950 7735 1971
rect 7801 1950 7831 1971
rect 7897 1950 7927 1971
rect 7993 1950 8023 1971
rect 8089 1950 8119 1971
rect 8185 1950 8215 1971
rect 8281 1950 8311 1971
rect 8377 1950 8407 1971
rect 8473 1950 8503 1971
rect 8569 1950 8599 1971
rect 8665 1950 8695 1971
rect 8761 1950 8791 1971
rect 8857 1950 8887 1971
rect 8953 1950 8983 1971
rect 9049 1950 9079 1971
rect 9145 1950 9175 1971
rect 9241 1950 9271 1971
rect 9337 1950 9367 1971
rect 9422 1969 9463 1971
rect 9433 1950 9463 1969
rect 9529 1950 9559 1971
rect -1407 -2019 -1377 -2000
rect -1311 -2019 -1281 -2000
rect -1215 -2019 -1185 -2000
rect -1119 -2019 -1089 -2000
rect -1023 -2019 -993 -2000
rect -927 -2019 -897 -2000
rect -831 -2019 -801 -2000
rect -735 -2019 -705 -2000
rect -639 -2019 -609 -2000
rect -543 -2019 -513 -2000
rect -447 -2019 -417 -2000
rect -351 -2019 -321 -2000
rect -255 -2019 -225 -2000
rect -159 -2019 -129 -2000
rect -63 -2019 -33 -2000
rect 33 -2019 63 -2000
rect 129 -2019 159 -2000
rect 225 -2019 255 -2000
rect 321 -2019 351 -2000
rect 417 -2019 447 -2000
rect 513 -2019 543 -2000
rect 609 -2019 639 -2000
rect 705 -2019 735 -2000
rect 801 -2019 831 -2000
rect 897 -2019 927 -2000
rect 993 -2019 1023 -2000
rect 1089 -2019 1119 -2000
rect 1185 -2019 1215 -2000
rect 1281 -2019 1311 -2000
rect 1377 -2019 1407 -2000
rect -1428 -2049 1444 -2019
rect 3865 -2069 3895 -2050
rect 3961 -2069 3991 -2050
rect 4057 -2069 4087 -2050
rect 4153 -2069 4183 -2050
rect 4249 -2069 4279 -2050
rect 4345 -2069 4375 -2050
rect 4441 -2069 4471 -2050
rect 4537 -2069 4567 -2050
rect 4633 -2069 4663 -2050
rect 4729 -2069 4759 -2050
rect 4825 -2069 4855 -2050
rect 4921 -2069 4951 -2050
rect 5017 -2069 5047 -2050
rect 5113 -2069 5143 -2050
rect 5209 -2069 5239 -2050
rect 5305 -2069 5335 -2050
rect 5401 -2069 5431 -2050
rect 5497 -2069 5527 -2050
rect 5593 -2069 5623 -2050
rect 5689 -2069 5719 -2050
rect 5785 -2069 5815 -2050
rect 5881 -2069 5911 -2050
rect 5977 -2069 6007 -2050
rect 6073 -2069 6103 -2050
rect 6169 -2069 6199 -2050
rect 6265 -2069 6295 -2050
rect 6361 -2069 6391 -2050
rect 6457 -2069 6487 -2050
rect 6553 -2069 6583 -2050
rect 6649 -2069 6679 -2050
rect 6745 -2069 6775 -2050
rect 6841 -2069 6871 -2050
rect 6937 -2069 6967 -2050
rect 7033 -2069 7063 -2050
rect 7129 -2069 7159 -2050
rect 7225 -2069 7255 -2050
rect 7321 -2069 7351 -2050
rect 7417 -2069 7447 -2050
rect 7513 -2069 7543 -2050
rect 7609 -2069 7639 -2050
rect 7705 -2069 7735 -2050
rect 7801 -2069 7831 -2050
rect 7897 -2069 7927 -2050
rect 7993 -2069 8023 -2050
rect 8089 -2069 8119 -2050
rect 8185 -2069 8215 -2050
rect 8281 -2069 8311 -2050
rect 8377 -2069 8407 -2050
rect 8473 -2069 8503 -2050
rect 8569 -2069 8599 -2050
rect 8665 -2069 8695 -2050
rect 8761 -2069 8791 -2050
rect 8857 -2069 8887 -2050
rect 8953 -2069 8983 -2050
rect 9049 -2069 9079 -2050
rect 9145 -2069 9175 -2050
rect 9241 -2069 9271 -2050
rect 9337 -2069 9367 -2050
rect 9433 -2069 9463 -2050
rect 9529 -2069 9559 -2050
rect 3844 -2099 9596 -2069
<< polycont >>
rect -1572 2003 -1510 2071
rect 3696 1959 3756 2017
<< locali >>
rect -1584 2071 -1494 2087
rect -1584 2055 -1572 2071
rect -1608 2021 -1572 2055
rect -1584 2003 -1572 2021
rect -1510 2003 -1494 2071
rect 3684 2017 3778 2037
rect 3684 2005 3696 2017
rect -1584 1987 -1494 2003
rect -1457 1988 -1423 2004
rect -1457 -2004 -1423 -1988
rect -1361 1988 -1327 2004
rect -1361 -1999 -1327 -1988
rect -1265 1988 -1231 2004
rect -1362 -2051 -1326 -1999
rect -1265 -2004 -1231 -1988
rect -1169 1988 -1135 2004
rect -1169 -1999 -1135 -1988
rect -1073 1988 -1039 2004
rect -1170 -2051 -1134 -1999
rect -1073 -2004 -1039 -1988
rect -977 1988 -943 2004
rect -977 -1999 -943 -1988
rect -881 1988 -847 2004
rect -978 -2051 -942 -1999
rect -881 -2004 -847 -1988
rect -785 1988 -751 2004
rect -785 -1999 -751 -1988
rect -689 1988 -655 2004
rect -786 -2051 -750 -1999
rect -689 -2004 -655 -1988
rect -593 1988 -559 2004
rect -593 -1999 -559 -1988
rect -497 1988 -463 2004
rect -594 -2051 -558 -1999
rect -497 -2004 -463 -1988
rect -401 1988 -367 2004
rect -401 -1999 -367 -1988
rect -305 1988 -271 2004
rect -402 -2051 -366 -1999
rect -305 -2004 -271 -1988
rect -209 1988 -175 2004
rect -209 -1999 -175 -1988
rect -113 1988 -79 2004
rect -210 -2051 -174 -1999
rect -113 -2004 -79 -1988
rect -17 1988 17 2004
rect -17 -1999 17 -1988
rect 79 1988 113 2004
rect -18 -2051 18 -1999
rect 79 -2004 113 -1988
rect 175 1988 209 2004
rect 175 -1999 209 -1988
rect 271 1988 305 2004
rect 174 -2051 210 -1999
rect 271 -2004 305 -1988
rect 367 1988 401 2004
rect 367 -1999 401 -1988
rect 463 1988 497 2004
rect 366 -2051 402 -1999
rect 463 -2004 497 -1988
rect 559 1988 593 2004
rect 559 -1999 593 -1988
rect 655 1988 689 2004
rect 558 -2051 594 -1999
rect 655 -2004 689 -1988
rect 751 1988 785 2004
rect 751 -1999 785 -1988
rect 847 1988 881 2004
rect 750 -2051 786 -1999
rect 847 -2004 881 -1988
rect 943 1988 977 2004
rect 943 -1999 977 -1988
rect 1039 1988 1073 2004
rect 942 -2051 978 -1999
rect 1039 -2004 1073 -1988
rect 1135 1988 1169 2004
rect 1135 -1999 1169 -1988
rect 1231 1988 1265 2004
rect 1134 -2051 1170 -1999
rect 1231 -2004 1265 -1988
rect 1327 1988 1361 2004
rect 1327 -1999 1361 -1988
rect 1423 1988 1457 2004
rect 3664 1971 3696 2005
rect 3684 1959 3696 1971
rect 3756 1959 3778 2017
rect 3684 1937 3778 1959
rect 3815 1938 3849 1954
rect 1326 -2051 1362 -1999
rect 1423 -2004 1457 -1988
rect -1418 -2061 1414 -2051
rect 3815 -2054 3849 -2038
rect 3911 1938 3945 1954
rect 3911 -2049 3945 -2038
rect 4007 1938 4041 1954
rect -1418 -2097 -1400 -2061
rect 1394 -2097 1414 -2061
rect -1418 -2105 1414 -2097
rect 3910 -2101 3946 -2049
rect 4007 -2054 4041 -2038
rect 4103 1938 4137 1954
rect 4103 -2049 4137 -2038
rect 4199 1938 4233 1954
rect 4102 -2101 4138 -2049
rect 4199 -2054 4233 -2038
rect 4295 1938 4329 1954
rect 4295 -2049 4329 -2038
rect 4391 1938 4425 1954
rect 4294 -2101 4330 -2049
rect 4391 -2054 4425 -2038
rect 4487 1938 4521 1954
rect 4487 -2049 4521 -2038
rect 4583 1938 4617 1954
rect 4486 -2101 4522 -2049
rect 4583 -2054 4617 -2038
rect 4679 1938 4713 1954
rect 4679 -2049 4713 -2038
rect 4775 1938 4809 1954
rect 4678 -2101 4714 -2049
rect 4775 -2054 4809 -2038
rect 4871 1938 4905 1954
rect 4871 -2049 4905 -2038
rect 4967 1938 5001 1954
rect 4870 -2101 4906 -2049
rect 4967 -2054 5001 -2038
rect 5063 1938 5097 1954
rect 5063 -2049 5097 -2038
rect 5159 1938 5193 1954
rect 5062 -2101 5098 -2049
rect 5159 -2054 5193 -2038
rect 5255 1938 5289 1954
rect 5255 -2049 5289 -2038
rect 5351 1938 5385 1954
rect 5254 -2101 5290 -2049
rect 5351 -2054 5385 -2038
rect 5447 1938 5481 1954
rect 5447 -2049 5481 -2038
rect 5543 1938 5577 1954
rect 5446 -2101 5482 -2049
rect 5543 -2054 5577 -2038
rect 5639 1938 5673 1954
rect 5639 -2049 5673 -2038
rect 5735 1938 5769 1954
rect 5638 -2101 5674 -2049
rect 5735 -2054 5769 -2038
rect 5831 1938 5865 1954
rect 5831 -2049 5865 -2038
rect 5927 1938 5961 1954
rect 5830 -2101 5866 -2049
rect 5927 -2054 5961 -2038
rect 6023 1938 6057 1954
rect 6023 -2049 6057 -2038
rect 6119 1938 6153 1954
rect 6022 -2101 6058 -2049
rect 6119 -2054 6153 -2038
rect 6215 1938 6249 1954
rect 6215 -2049 6249 -2038
rect 6311 1938 6345 1954
rect 6214 -2101 6250 -2049
rect 6311 -2054 6345 -2038
rect 6407 1938 6441 1954
rect 6407 -2049 6441 -2038
rect 6503 1938 6537 1954
rect 6406 -2101 6442 -2049
rect 6503 -2054 6537 -2038
rect 6599 1938 6633 1954
rect 6599 -2049 6633 -2038
rect 6695 1938 6729 1954
rect 6598 -2101 6634 -2049
rect 6695 -2054 6729 -2038
rect 6791 1938 6825 1954
rect 6791 -2049 6825 -2038
rect 6887 1938 6921 1954
rect 6790 -2101 6826 -2049
rect 6887 -2054 6921 -2038
rect 6983 1938 7017 1954
rect 6983 -2049 7017 -2038
rect 7079 1938 7113 1954
rect 6982 -2101 7018 -2049
rect 7079 -2054 7113 -2038
rect 7175 1938 7209 1954
rect 7175 -2049 7209 -2038
rect 7271 1938 7305 1954
rect 7174 -2101 7210 -2049
rect 7271 -2054 7305 -2038
rect 7367 1938 7401 1954
rect 7367 -2049 7401 -2038
rect 7463 1938 7497 1954
rect 7366 -2101 7402 -2049
rect 7463 -2054 7497 -2038
rect 7559 1938 7593 1954
rect 7559 -2049 7593 -2038
rect 7655 1938 7689 1954
rect 7558 -2101 7594 -2049
rect 7655 -2054 7689 -2038
rect 7751 1938 7785 1954
rect 7751 -2049 7785 -2038
rect 7847 1938 7881 1954
rect 7750 -2101 7786 -2049
rect 7847 -2054 7881 -2038
rect 7943 1938 7977 1954
rect 7943 -2049 7977 -2038
rect 8039 1938 8073 1954
rect 7942 -2101 7978 -2049
rect 8039 -2054 8073 -2038
rect 8135 1938 8169 1954
rect 8135 -2049 8169 -2038
rect 8231 1938 8265 1954
rect 8134 -2101 8170 -2049
rect 8231 -2054 8265 -2038
rect 8327 1938 8361 1954
rect 8327 -2049 8361 -2038
rect 8423 1938 8457 1954
rect 8326 -2101 8362 -2049
rect 8423 -2054 8457 -2038
rect 8519 1938 8553 1954
rect 8519 -2049 8553 -2038
rect 8615 1938 8649 1954
rect 8518 -2101 8554 -2049
rect 8615 -2054 8649 -2038
rect 8711 1938 8745 1954
rect 8711 -2049 8745 -2038
rect 8807 1938 8841 1954
rect 8710 -2101 8746 -2049
rect 8807 -2054 8841 -2038
rect 8903 1938 8937 1954
rect 8903 -2049 8937 -2038
rect 8999 1938 9033 1954
rect 8902 -2101 8938 -2049
rect 8999 -2054 9033 -2038
rect 9095 1938 9129 1954
rect 9095 -2049 9129 -2038
rect 9191 1938 9225 1954
rect 9094 -2101 9130 -2049
rect 9191 -2054 9225 -2038
rect 9287 1938 9321 1954
rect 9287 -2049 9321 -2038
rect 9383 1938 9417 1954
rect 9286 -2101 9322 -2049
rect 9383 -2054 9417 -2038
rect 9479 1938 9513 1954
rect 9479 -2049 9513 -2038
rect 9575 1938 9609 1954
rect 9478 -2101 9514 -2049
rect 9575 -2054 9609 -2038
rect -1362 -2140 -1326 -2105
rect -1170 -2140 -1134 -2105
rect -978 -2140 -942 -2105
rect -786 -2140 -750 -2105
rect -594 -2140 -558 -2105
rect -402 -2140 -366 -2105
rect -210 -2140 -174 -2105
rect -18 -2140 18 -2105
rect 174 -2140 210 -2105
rect 366 -2140 402 -2105
rect 558 -2140 594 -2105
rect 750 -2140 786 -2105
rect 942 -2140 978 -2105
rect 1134 -2140 1170 -2105
rect 1326 -2140 1362 -2105
rect 3860 -2111 9566 -2101
rect -1537 -2174 -1473 -2140
rect 1477 -2174 1534 -2140
rect 3860 -2147 3872 -2111
rect 6666 -2147 6752 -2111
rect 9546 -2147 9566 -2111
rect 3860 -2155 9566 -2147
rect 3910 -2190 3946 -2155
rect 4102 -2190 4138 -2155
rect 4294 -2190 4330 -2155
rect 4486 -2190 4522 -2155
rect 4678 -2190 4714 -2155
rect 4870 -2190 4906 -2155
rect 5062 -2190 5098 -2155
rect 5254 -2190 5290 -2155
rect 5446 -2190 5482 -2155
rect 5638 -2190 5674 -2155
rect 5830 -2190 5866 -2155
rect 6022 -2190 6058 -2155
rect 6214 -2190 6250 -2155
rect 6406 -2190 6442 -2155
rect 6598 -2190 6634 -2155
rect 6790 -2190 6826 -2155
rect 6982 -2190 7018 -2155
rect 7174 -2190 7210 -2155
rect 7366 -2190 7402 -2155
rect 7558 -2190 7594 -2155
rect 7750 -2190 7786 -2155
rect 7942 -2190 7978 -2155
rect 8134 -2190 8170 -2155
rect 8326 -2190 8362 -2155
rect 8518 -2190 8554 -2155
rect 8710 -2190 8746 -2155
rect 8902 -2190 8938 -2155
rect 9094 -2190 9130 -2155
rect 9286 -2190 9322 -2155
rect 9478 -2190 9514 -2155
rect 3735 -2224 3799 -2190
rect 9629 -2224 9686 -2190
<< viali >>
rect -1457 -1988 -1423 1988
rect -1361 -1988 -1327 1988
rect -1265 -1988 -1231 1988
rect -1169 -1988 -1135 1988
rect -1073 -1988 -1039 1988
rect -977 -1988 -943 1988
rect -881 -1988 -847 1988
rect -785 -1988 -751 1988
rect -689 -1988 -655 1988
rect -593 -1988 -559 1988
rect -497 -1988 -463 1988
rect -401 -1988 -367 1988
rect -305 -1988 -271 1988
rect -209 -1988 -175 1988
rect -113 -1988 -79 1988
rect -17 -1988 17 1988
rect 79 -1988 113 1988
rect 175 -1988 209 1988
rect 271 -1988 305 1988
rect 367 -1988 401 1988
rect 463 -1988 497 1988
rect 559 -1988 593 1988
rect 655 -1988 689 1988
rect 751 -1988 785 1988
rect 847 -1988 881 1988
rect 943 -1988 977 1988
rect 1039 -1988 1073 1988
rect 1135 -1988 1169 1988
rect 1231 -1988 1265 1988
rect 1327 -1988 1361 1988
rect 1423 -1988 1457 1988
rect 3700 1961 3752 2015
rect 3815 -2038 3849 1938
rect 3911 -2038 3945 1938
rect 4007 -2038 4041 1938
rect -1400 -2097 1394 -2061
rect 4103 -2038 4137 1938
rect 4199 -2038 4233 1938
rect 4295 -2038 4329 1938
rect 4391 -2038 4425 1938
rect 4487 -2038 4521 1938
rect 4583 -2038 4617 1938
rect 4679 -2038 4713 1938
rect 4775 -2038 4809 1938
rect 4871 -2038 4905 1938
rect 4967 -2038 5001 1938
rect 5063 -2038 5097 1938
rect 5159 -2038 5193 1938
rect 5255 -2038 5289 1938
rect 5351 -2038 5385 1938
rect 5447 -2038 5481 1938
rect 5543 -2038 5577 1938
rect 5639 -2038 5673 1938
rect 5735 -2038 5769 1938
rect 5831 -2038 5865 1938
rect 5927 -2038 5961 1938
rect 6023 -2038 6057 1938
rect 6119 -2038 6153 1938
rect 6215 -2038 6249 1938
rect 6311 -2038 6345 1938
rect 6407 -2038 6441 1938
rect 6503 -2038 6537 1938
rect 6599 -2038 6633 1938
rect 6695 -2038 6729 1938
rect 6791 -2038 6825 1938
rect 6887 -2038 6921 1938
rect 6983 -2038 7017 1938
rect 7079 -2038 7113 1938
rect 7175 -2038 7209 1938
rect 7271 -2038 7305 1938
rect 7367 -2038 7401 1938
rect 7463 -2038 7497 1938
rect 7559 -2038 7593 1938
rect 7655 -2038 7689 1938
rect 7751 -2038 7785 1938
rect 7847 -2038 7881 1938
rect 7943 -2038 7977 1938
rect 8039 -2038 8073 1938
rect 8135 -2038 8169 1938
rect 8231 -2038 8265 1938
rect 8327 -2038 8361 1938
rect 8423 -2038 8457 1938
rect 8519 -2038 8553 1938
rect 8615 -2038 8649 1938
rect 8711 -2038 8745 1938
rect 8807 -2038 8841 1938
rect 8903 -2038 8937 1938
rect 8999 -2038 9033 1938
rect 9095 -2038 9129 1938
rect 9191 -2038 9225 1938
rect 9287 -2038 9321 1938
rect 9383 -2038 9417 1938
rect 9479 -2038 9513 1938
rect 9575 -2038 9609 1938
rect 3872 -2147 6666 -2111
rect 6752 -2147 9546 -2111
<< metal1 >>
rect -116 2543 5194 2603
rect -116 2159 -74 2543
rect 5156 2161 5194 2543
rect -1472 2115 1462 2159
rect -1462 2000 -1418 2115
rect -1270 2000 -1226 2115
rect -1078 2000 -1034 2115
rect -1463 1988 -1417 2000
rect -1463 -1988 -1457 1988
rect -1423 -1988 -1417 1988
rect -1463 -2000 -1417 -1988
rect -1367 1988 -1321 2000
rect -1367 -1988 -1361 1988
rect -1327 -1988 -1321 1988
rect -1367 -2000 -1321 -1988
rect -1271 1988 -1225 2000
rect -1271 -1988 -1265 1988
rect -1231 -1988 -1225 1988
rect -1271 -2000 -1225 -1988
rect -1175 1988 -1129 2000
rect -1175 -1988 -1169 1988
rect -1135 -1988 -1129 1988
rect -1175 -2000 -1129 -1988
rect -1079 1999 -1034 2000
rect -1079 1988 -1033 1999
rect -1079 -1988 -1073 1988
rect -1039 -1988 -1033 1988
rect -1079 -2000 -1033 -1988
rect -983 1988 -937 2000
rect -886 1999 -842 2115
rect -983 -1988 -977 1988
rect -943 -1988 -937 1988
rect -983 -2000 -937 -1988
rect -887 1988 -841 1999
rect -887 -1988 -881 1988
rect -847 -1988 -841 1988
rect -887 -2000 -841 -1988
rect -791 1988 -745 2000
rect -694 1999 -650 2115
rect -502 2000 -458 2115
rect -310 2000 -266 2115
rect -118 2000 -74 2115
rect 74 2001 118 2115
rect 74 2000 119 2001
rect -791 -1988 -785 1988
rect -751 -1988 -745 1988
rect -791 -2000 -745 -1988
rect -695 1988 -649 1999
rect -695 -1988 -689 1988
rect -655 -1988 -649 1988
rect -695 -2000 -649 -1988
rect -599 1988 -553 2000
rect -502 1999 -457 2000
rect -599 -1988 -593 1988
rect -559 -1988 -553 1988
rect -599 -2000 -553 -1988
rect -503 1988 -457 1999
rect -503 -1988 -497 1988
rect -463 -1988 -457 1988
rect -503 -2000 -457 -1988
rect -407 1988 -361 2000
rect -407 -1988 -401 1988
rect -367 -1988 -361 1988
rect -407 -2000 -361 -1988
rect -311 1988 -265 2000
rect -311 -1988 -305 1988
rect -271 -1988 -265 1988
rect -311 -2000 -265 -1988
rect -215 1988 -169 2000
rect -215 -1988 -209 1988
rect -175 -1988 -169 1988
rect -215 -1999 -169 -1988
rect -119 1988 -73 2000
rect -119 -1988 -113 1988
rect -79 -1988 -73 1988
rect -215 -2000 -174 -1999
rect -119 -2000 -73 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 73 1988 119 2000
rect 73 -1988 79 1988
rect 113 -1988 119 1988
rect 73 -2000 119 -1988
rect 169 1988 215 2000
rect 266 1999 310 2115
rect 458 2000 502 2115
rect 650 2000 694 2115
rect 842 2000 886 2115
rect 1034 2000 1078 2115
rect 1226 2000 1270 2115
rect 1418 2000 1462 2115
rect 5156 2109 5198 2161
rect 8036 2109 8078 2161
rect 3800 2065 9614 2109
rect 169 -1988 175 1988
rect 209 -1988 215 1988
rect 169 -2000 215 -1988
rect 265 1988 311 1999
rect 265 -1988 271 1988
rect 305 -1988 311 1988
rect 265 -2000 311 -1988
rect 361 1988 407 2000
rect 361 -1988 367 1988
rect 401 -1988 407 1988
rect 361 -2000 407 -1988
rect 457 1999 502 2000
rect 457 1988 503 1999
rect 457 -1988 463 1988
rect 497 -1988 503 1988
rect 457 -2000 503 -1988
rect 553 1988 599 2000
rect 650 1999 695 2000
rect 553 -1988 559 1988
rect 593 -1988 599 1988
rect 553 -2000 599 -1988
rect 649 1988 695 1999
rect 649 -1988 655 1988
rect 689 -1988 695 1988
rect 649 -2000 695 -1988
rect 745 1988 791 2000
rect 842 1999 887 2000
rect 745 -1988 751 1988
rect 785 -1988 791 1988
rect 745 -2000 791 -1988
rect 841 1988 887 1999
rect 841 -1988 847 1988
rect 881 -1988 887 1988
rect 841 -2000 887 -1988
rect 937 1988 983 2000
rect 1034 1999 1079 2000
rect 937 -1988 943 1988
rect 977 -1988 983 1988
rect 937 -2000 983 -1988
rect 1033 1988 1079 1999
rect 1033 -1988 1039 1988
rect 1073 -1988 1079 1988
rect 1033 -2000 1079 -1988
rect 1129 1988 1175 2000
rect 1129 -1988 1135 1988
rect 1169 -1988 1175 1988
rect 1129 -2000 1175 -1988
rect 1225 1999 1270 2000
rect 1225 1988 1271 1999
rect 1225 -1988 1231 1988
rect 1265 -1988 1271 1988
rect 1225 -2000 1271 -1988
rect 1321 1988 1367 2000
rect 1321 -1988 1327 1988
rect 1361 -1988 1367 1988
rect 1321 -1999 1367 -1988
rect 1417 1999 1462 2000
rect 3692 2015 3762 2031
rect 1417 1988 1463 1999
rect 1417 -1988 1423 1988
rect 1457 -1988 1463 1988
rect 1321 -2000 1362 -1999
rect 1417 -2000 1463 -1988
rect 3692 1961 3700 2015
rect 3752 1961 3762 2015
rect -1418 -2061 1414 -2051
rect -1418 -2097 -1400 -2061
rect 1394 -2097 1414 -2061
rect -1418 -2105 1414 -2097
rect 3692 -2101 3762 1961
rect 3810 1950 3854 2065
rect 4002 1950 4046 2065
rect 4194 1950 4238 2065
rect 3809 1938 3855 1950
rect 3809 -2038 3815 1938
rect 3849 -2038 3855 1938
rect 3809 -2050 3855 -2038
rect 3905 1938 3951 1950
rect 3905 -2038 3911 1938
rect 3945 -2038 3951 1938
rect 3905 -2050 3951 -2038
rect 4001 1938 4047 1950
rect 4001 -2038 4007 1938
rect 4041 -2038 4047 1938
rect 4001 -2050 4047 -2038
rect 4097 1938 4143 1950
rect 4097 -2038 4103 1938
rect 4137 -2038 4143 1938
rect 4097 -2050 4143 -2038
rect 4193 1949 4238 1950
rect 4193 1938 4239 1949
rect 4193 -2038 4199 1938
rect 4233 -2038 4239 1938
rect 4193 -2050 4239 -2038
rect 4289 1938 4335 1950
rect 4386 1949 4430 2065
rect 4289 -2038 4295 1938
rect 4329 -2038 4335 1938
rect 4289 -2050 4335 -2038
rect 4385 1938 4431 1949
rect 4385 -2038 4391 1938
rect 4425 -2038 4431 1938
rect 4385 -2050 4431 -2038
rect 4481 1938 4527 1950
rect 4578 1949 4622 2065
rect 4770 1950 4814 2065
rect 4962 1950 5006 2065
rect 5154 1950 5198 2065
rect 5346 1951 5390 2065
rect 5346 1950 5391 1951
rect 4481 -2038 4487 1938
rect 4521 -2038 4527 1938
rect 4481 -2050 4527 -2038
rect 4577 1938 4623 1949
rect 4577 -2038 4583 1938
rect 4617 -2038 4623 1938
rect 4577 -2050 4623 -2038
rect 4673 1938 4719 1950
rect 4770 1949 4815 1950
rect 4673 -2038 4679 1938
rect 4713 -2038 4719 1938
rect 4673 -2050 4719 -2038
rect 4769 1938 4815 1949
rect 4769 -2038 4775 1938
rect 4809 -2038 4815 1938
rect 4769 -2050 4815 -2038
rect 4865 1938 4911 1950
rect 4865 -2038 4871 1938
rect 4905 -2038 4911 1938
rect 4865 -2050 4911 -2038
rect 4961 1938 5007 1950
rect 4961 -2038 4967 1938
rect 5001 -2038 5007 1938
rect 4961 -2050 5007 -2038
rect 5057 1938 5103 1950
rect 5057 -2038 5063 1938
rect 5097 -2038 5103 1938
rect 5057 -2049 5103 -2038
rect 5153 1938 5199 1950
rect 5153 -2038 5159 1938
rect 5193 -2038 5199 1938
rect 5057 -2050 5098 -2049
rect 5153 -2050 5199 -2038
rect 5249 1938 5295 1950
rect 5249 -2038 5255 1938
rect 5289 -2038 5295 1938
rect 5249 -2050 5295 -2038
rect 5345 1938 5391 1950
rect 5345 -2038 5351 1938
rect 5385 -2038 5391 1938
rect 5345 -2050 5391 -2038
rect 5441 1938 5487 1950
rect 5538 1949 5582 2065
rect 5730 1950 5774 2065
rect 5922 1950 5966 2065
rect 6114 1950 6158 2065
rect 6306 1950 6350 2065
rect 6498 1950 6542 2065
rect 6690 1950 6734 2065
rect 6882 1950 6926 2065
rect 7074 1950 7118 2065
rect 5441 -2038 5447 1938
rect 5481 -2038 5487 1938
rect 5441 -2050 5487 -2038
rect 5537 1938 5583 1949
rect 5537 -2038 5543 1938
rect 5577 -2038 5583 1938
rect 5537 -2050 5583 -2038
rect 5633 1938 5679 1950
rect 5633 -2038 5639 1938
rect 5673 -2038 5679 1938
rect 5633 -2050 5679 -2038
rect 5729 1949 5774 1950
rect 5729 1938 5775 1949
rect 5729 -2038 5735 1938
rect 5769 -2038 5775 1938
rect 5729 -2050 5775 -2038
rect 5825 1938 5871 1950
rect 5922 1949 5967 1950
rect 5825 -2038 5831 1938
rect 5865 -2038 5871 1938
rect 5825 -2050 5871 -2038
rect 5921 1938 5967 1949
rect 5921 -2038 5927 1938
rect 5961 -2038 5967 1938
rect 5921 -2050 5967 -2038
rect 6017 1938 6063 1950
rect 6114 1949 6159 1950
rect 6017 -2038 6023 1938
rect 6057 -2038 6063 1938
rect 6017 -2050 6063 -2038
rect 6113 1938 6159 1949
rect 6113 -2038 6119 1938
rect 6153 -2038 6159 1938
rect 6113 -2050 6159 -2038
rect 6209 1938 6255 1950
rect 6306 1949 6351 1950
rect 6209 -2038 6215 1938
rect 6249 -2038 6255 1938
rect 6209 -2050 6255 -2038
rect 6305 1938 6351 1949
rect 6305 -2038 6311 1938
rect 6345 -2038 6351 1938
rect 6305 -2050 6351 -2038
rect 6401 1938 6447 1950
rect 6401 -2038 6407 1938
rect 6441 -2038 6447 1938
rect 6401 -2050 6447 -2038
rect 6497 1949 6542 1950
rect 6497 1938 6543 1949
rect 6497 -2038 6503 1938
rect 6537 -2038 6543 1938
rect 6497 -2050 6543 -2038
rect 6593 1938 6639 1950
rect 6593 -2038 6599 1938
rect 6633 -2038 6639 1938
rect 6593 -2049 6639 -2038
rect 6689 1949 6734 1950
rect 6689 1938 6735 1949
rect 6689 -2038 6695 1938
rect 6729 -2038 6735 1938
rect 6593 -2050 6634 -2049
rect 6689 -2050 6735 -2038
rect 6785 1938 6831 1950
rect 6785 -2038 6791 1938
rect 6825 -2038 6831 1938
rect 6785 -2050 6831 -2038
rect 6881 1938 6927 1950
rect 6881 -2038 6887 1938
rect 6921 -2038 6927 1938
rect 6881 -2050 6927 -2038
rect 6977 1938 7023 1950
rect 6977 -2038 6983 1938
rect 7017 -2038 7023 1938
rect 6977 -2050 7023 -2038
rect 7073 1949 7118 1950
rect 7073 1938 7119 1949
rect 7073 -2038 7079 1938
rect 7113 -2038 7119 1938
rect 7073 -2050 7119 -2038
rect 7169 1938 7215 1950
rect 7266 1949 7310 2065
rect 7169 -2038 7175 1938
rect 7209 -2038 7215 1938
rect 7169 -2050 7215 -2038
rect 7265 1938 7311 1949
rect 7265 -2038 7271 1938
rect 7305 -2038 7311 1938
rect 7265 -2050 7311 -2038
rect 7361 1938 7407 1950
rect 7458 1949 7502 2065
rect 7650 1950 7694 2065
rect 7842 1950 7886 2065
rect 8034 1950 8078 2065
rect 8226 1951 8270 2065
rect 8226 1950 8271 1951
rect 7361 -2038 7367 1938
rect 7401 -2038 7407 1938
rect 7361 -2050 7407 -2038
rect 7457 1938 7503 1949
rect 7457 -2038 7463 1938
rect 7497 -2038 7503 1938
rect 7457 -2050 7503 -2038
rect 7553 1938 7599 1950
rect 7650 1949 7695 1950
rect 7553 -2038 7559 1938
rect 7593 -2038 7599 1938
rect 7553 -2050 7599 -2038
rect 7649 1938 7695 1949
rect 7649 -2038 7655 1938
rect 7689 -2038 7695 1938
rect 7649 -2050 7695 -2038
rect 7745 1938 7791 1950
rect 7745 -2038 7751 1938
rect 7785 -2038 7791 1938
rect 7745 -2050 7791 -2038
rect 7841 1938 7887 1950
rect 7841 -2038 7847 1938
rect 7881 -2038 7887 1938
rect 7841 -2050 7887 -2038
rect 7937 1938 7983 1950
rect 7937 -2038 7943 1938
rect 7977 -2038 7983 1938
rect 7937 -2049 7983 -2038
rect 8033 1938 8079 1950
rect 8033 -2038 8039 1938
rect 8073 -2038 8079 1938
rect 7937 -2050 7978 -2049
rect 8033 -2050 8079 -2038
rect 8129 1938 8175 1950
rect 8129 -2038 8135 1938
rect 8169 -2038 8175 1938
rect 8129 -2050 8175 -2038
rect 8225 1938 8271 1950
rect 8225 -2038 8231 1938
rect 8265 -2038 8271 1938
rect 8225 -2050 8271 -2038
rect 8321 1938 8367 1950
rect 8418 1949 8462 2065
rect 8610 1950 8654 2065
rect 8802 1950 8846 2065
rect 8994 1950 9038 2065
rect 9186 1950 9230 2065
rect 9378 1950 9422 2065
rect 9570 1950 9614 2065
rect 8321 -2038 8327 1938
rect 8361 -2038 8367 1938
rect 8321 -2050 8367 -2038
rect 8417 1938 8463 1949
rect 8417 -2038 8423 1938
rect 8457 -2038 8463 1938
rect 8417 -2050 8463 -2038
rect 8513 1938 8559 1950
rect 8513 -2038 8519 1938
rect 8553 -2038 8559 1938
rect 8513 -2050 8559 -2038
rect 8609 1949 8654 1950
rect 8609 1938 8655 1949
rect 8609 -2038 8615 1938
rect 8649 -2038 8655 1938
rect 8609 -2050 8655 -2038
rect 8705 1938 8751 1950
rect 8802 1949 8847 1950
rect 8705 -2038 8711 1938
rect 8745 -2038 8751 1938
rect 8705 -2050 8751 -2038
rect 8801 1938 8847 1949
rect 8801 -2038 8807 1938
rect 8841 -2038 8847 1938
rect 8801 -2050 8847 -2038
rect 8897 1938 8943 1950
rect 8994 1949 9039 1950
rect 8897 -2038 8903 1938
rect 8937 -2038 8943 1938
rect 8897 -2050 8943 -2038
rect 8993 1938 9039 1949
rect 8993 -2038 8999 1938
rect 9033 -2038 9039 1938
rect 8993 -2050 9039 -2038
rect 9089 1938 9135 1950
rect 9186 1949 9231 1950
rect 9089 -2038 9095 1938
rect 9129 -2038 9135 1938
rect 9089 -2050 9135 -2038
rect 9185 1938 9231 1949
rect 9185 -2038 9191 1938
rect 9225 -2038 9231 1938
rect 9185 -2050 9231 -2038
rect 9281 1938 9327 1950
rect 9281 -2038 9287 1938
rect 9321 -2038 9327 1938
rect 9281 -2050 9327 -2038
rect 9377 1949 9422 1950
rect 9377 1938 9423 1949
rect 9377 -2038 9383 1938
rect 9417 -2038 9423 1938
rect 9377 -2050 9423 -2038
rect 9473 1938 9519 1950
rect 9473 -2038 9479 1938
rect 9513 -2038 9519 1938
rect 9473 -2049 9519 -2038
rect 9569 1949 9614 1950
rect 9569 1938 9615 1949
rect 9569 -2038 9575 1938
rect 9609 -2038 9615 1938
rect 9473 -2050 9514 -2049
rect 9569 -2050 9615 -2038
rect -20 -2213 18 -2105
rect 3692 -2111 9566 -2101
rect 3692 -2147 3872 -2111
rect 6666 -2147 6752 -2111
rect 9546 -2147 9566 -2111
rect 3692 -2155 9566 -2147
rect 5252 -2263 5290 -2155
rect 8132 -2345 8170 -2155
<< labels >>
rlabel locali -1608 2039 -1608 2039 7 CKS
rlabel metal1 -94 2603 -94 2603 1 VX
rlabel metal1 -2 -2213 -2 -2213 5 VN
rlabel metal1 8150 -2345 8150 -2345 5 OUT
<< properties >>
string FIXED_BBOX -1554 -2157 1554 2157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20 l 0.150 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
