magic
tech sky130A
magscale 1 2
timestamp 1661709240
<< checkpaint >>
rect -1313 2276 6341 2329
rect -1313 2255 11422 2276
rect -1313 -713 14583 2255
rect 3768 -766 14583 -713
rect 8849 -819 14583 -766
<< error_p >>
rect 229 931 287 937
rect 421 931 479 937
rect 613 931 671 937
rect 805 931 863 937
rect 997 931 1055 937
rect 1189 931 1247 937
rect 1381 931 1439 937
rect 1573 931 1631 937
rect 1765 931 1823 937
rect 1957 931 2015 937
rect 2149 931 2207 937
rect 2341 931 2399 937
rect 2533 931 2591 937
rect 2725 931 2783 937
rect 2917 931 2975 937
rect 3109 931 3167 937
rect 3301 931 3359 937
rect 3493 931 3551 937
rect 3685 931 3743 937
rect 3877 931 3935 937
rect 4069 931 4127 937
rect 4261 931 4319 937
rect 4453 931 4511 937
rect 4645 931 4703 937
rect 4837 931 4895 937
rect 229 897 241 931
rect 421 897 433 931
rect 613 897 625 931
rect 805 897 817 931
rect 997 897 1009 931
rect 1189 897 1201 931
rect 1381 897 1393 931
rect 1573 897 1585 931
rect 1765 897 1777 931
rect 1957 897 1969 931
rect 2149 897 2161 931
rect 2341 897 2353 931
rect 2533 897 2545 931
rect 2725 897 2737 931
rect 2917 897 2929 931
rect 3109 897 3121 931
rect 3301 897 3313 931
rect 3493 897 3505 931
rect 3685 897 3697 931
rect 3877 897 3889 931
rect 4069 897 4081 931
rect 4261 897 4273 931
rect 4453 897 4465 931
rect 4645 897 4657 931
rect 4837 897 4849 931
rect 229 891 287 897
rect 421 891 479 897
rect 613 891 671 897
rect 805 891 863 897
rect 997 891 1055 897
rect 1189 891 1247 897
rect 1381 891 1439 897
rect 1573 891 1631 897
rect 1765 891 1823 897
rect 1957 891 2015 897
rect 2149 891 2207 897
rect 2341 891 2399 897
rect 2533 891 2591 897
rect 2725 891 2783 897
rect 2917 891 2975 897
rect 3109 891 3167 897
rect 3301 891 3359 897
rect 3493 891 3551 897
rect 3685 891 3743 897
rect 3877 891 3935 897
rect 4069 891 4127 897
rect 4261 891 4319 897
rect 4453 891 4511 897
rect 4645 891 4703 897
rect 4837 891 4895 897
rect 133 719 191 725
rect 325 719 383 725
rect 517 719 575 725
rect 709 719 767 725
rect 901 719 959 725
rect 1093 719 1151 725
rect 1285 719 1343 725
rect 1477 719 1535 725
rect 1669 719 1727 725
rect 1861 719 1919 725
rect 2053 719 2111 725
rect 2245 719 2303 725
rect 2437 719 2495 725
rect 2629 719 2687 725
rect 2821 719 2879 725
rect 3013 719 3071 725
rect 3205 719 3263 725
rect 3397 719 3455 725
rect 3589 719 3647 725
rect 3781 719 3839 725
rect 3973 719 4031 725
rect 4165 719 4223 725
rect 4357 719 4415 725
rect 4549 719 4607 725
rect 4741 719 4799 725
rect 133 685 145 719
rect 325 685 337 719
rect 517 685 529 719
rect 709 685 721 719
rect 901 685 913 719
rect 1093 685 1105 719
rect 1285 685 1297 719
rect 1477 685 1489 719
rect 1669 685 1681 719
rect 1861 685 1873 719
rect 2053 685 2065 719
rect 2245 685 2257 719
rect 2437 685 2449 719
rect 2629 685 2641 719
rect 2821 685 2833 719
rect 3013 685 3025 719
rect 3205 685 3217 719
rect 3397 685 3409 719
rect 3589 685 3601 719
rect 3781 685 3793 719
rect 3973 685 3985 719
rect 4165 685 4177 719
rect 4357 685 4369 719
rect 4549 685 4561 719
rect 4741 685 4753 719
rect 133 679 191 685
rect 325 679 383 685
rect 517 679 575 685
rect 709 679 767 685
rect 901 679 959 685
rect 1093 679 1151 685
rect 1285 679 1343 685
rect 1477 679 1535 685
rect 1669 679 1727 685
rect 1861 679 1919 685
rect 2053 679 2111 685
rect 2245 679 2303 685
rect 2437 679 2495 685
rect 2629 679 2687 685
rect 2821 679 2879 685
rect 3013 679 3071 685
rect 3205 679 3263 685
rect 3397 679 3455 685
rect 3589 679 3647 685
rect 3781 679 3839 685
rect 3973 679 4031 685
rect 4165 679 4223 685
rect 4357 679 4415 685
rect 4549 679 4607 685
rect 4741 679 4799 685
use sky130_fd_pr__pfet_01v8_2DBJRP  XM1
timestamp 0
transform 1 0 2514 0 1 808
box -2567 -261 2567 261
use sky130_fd_pr__pfet_01v8_2DBJRP  XM2
timestamp 0
transform 1 0 7595 0 1 755
box -2567 -261 2567 261
use sky130_fd_pr__nfet_01v8_ZEAV3T  XM3
timestamp 0
transform 1 0 11716 0 1 718
box -1607 -277 1607 277
<< end >>
