magic
tech sky130A
magscale 1 2
timestamp 1661696654
<< nmos >>
rect -2847 -1000 -2817 1000
rect -2751 -1000 -2721 1000
rect -2655 -1000 -2625 1000
rect -2559 -1000 -2529 1000
rect -2463 -1000 -2433 1000
rect -2367 -1000 -2337 1000
rect -2271 -1000 -2241 1000
rect -2175 -1000 -2145 1000
rect -2079 -1000 -2049 1000
rect -1983 -1000 -1953 1000
rect -1887 -1000 -1857 1000
rect -1791 -1000 -1761 1000
rect -1695 -1000 -1665 1000
rect -1599 -1000 -1569 1000
rect -1503 -1000 -1473 1000
rect -1407 -1000 -1377 1000
rect -1311 -1000 -1281 1000
rect -1215 -1000 -1185 1000
rect -1119 -1000 -1089 1000
rect -1023 -1000 -993 1000
rect -927 -1000 -897 1000
rect -831 -1000 -801 1000
rect -735 -1000 -705 1000
rect -639 -1000 -609 1000
rect -543 -1000 -513 1000
rect -447 -1000 -417 1000
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
rect 417 -1000 447 1000
rect 513 -1000 543 1000
rect 609 -1000 639 1000
rect 705 -1000 735 1000
rect 801 -1000 831 1000
rect 897 -1000 927 1000
rect 993 -1000 1023 1000
rect 1089 -1000 1119 1000
rect 1185 -1000 1215 1000
rect 1281 -1000 1311 1000
rect 1377 -1000 1407 1000
rect 1473 -1000 1503 1000
rect 1569 -1000 1599 1000
rect 1665 -1000 1695 1000
rect 1761 -1000 1791 1000
rect 1857 -1000 1887 1000
rect 1953 -1000 1983 1000
rect 2049 -1000 2079 1000
rect 2145 -1000 2175 1000
rect 2241 -1000 2271 1000
rect 2337 -1000 2367 1000
rect 2433 -1000 2463 1000
rect 2529 -1000 2559 1000
rect 2625 -1000 2655 1000
rect 2721 -1000 2751 1000
rect 2817 -1000 2847 1000
<< ndiff >>
rect -2909 988 -2847 1000
rect -2909 -988 -2897 988
rect -2863 -988 -2847 988
rect -2909 -1000 -2847 -988
rect -2817 988 -2751 1000
rect -2817 -988 -2801 988
rect -2767 -988 -2751 988
rect -2817 -1000 -2751 -988
rect -2721 988 -2655 1000
rect -2721 -988 -2705 988
rect -2671 -988 -2655 988
rect -2721 -1000 -2655 -988
rect -2625 988 -2559 1000
rect -2625 -988 -2609 988
rect -2575 -988 -2559 988
rect -2625 -1000 -2559 -988
rect -2529 988 -2463 1000
rect -2529 -988 -2513 988
rect -2479 -988 -2463 988
rect -2529 -1000 -2463 -988
rect -2433 988 -2367 1000
rect -2433 -988 -2417 988
rect -2383 -988 -2367 988
rect -2433 -1000 -2367 -988
rect -2337 988 -2271 1000
rect -2337 -988 -2321 988
rect -2287 -988 -2271 988
rect -2337 -1000 -2271 -988
rect -2241 988 -2175 1000
rect -2241 -988 -2225 988
rect -2191 -988 -2175 988
rect -2241 -1000 -2175 -988
rect -2145 988 -2079 1000
rect -2145 -988 -2129 988
rect -2095 -988 -2079 988
rect -2145 -1000 -2079 -988
rect -2049 988 -1983 1000
rect -2049 -988 -2033 988
rect -1999 -988 -1983 988
rect -2049 -1000 -1983 -988
rect -1953 988 -1887 1000
rect -1953 -988 -1937 988
rect -1903 -988 -1887 988
rect -1953 -1000 -1887 -988
rect -1857 988 -1791 1000
rect -1857 -988 -1841 988
rect -1807 -988 -1791 988
rect -1857 -1000 -1791 -988
rect -1761 988 -1695 1000
rect -1761 -988 -1745 988
rect -1711 -988 -1695 988
rect -1761 -1000 -1695 -988
rect -1665 988 -1599 1000
rect -1665 -988 -1649 988
rect -1615 -988 -1599 988
rect -1665 -1000 -1599 -988
rect -1569 988 -1503 1000
rect -1569 -988 -1553 988
rect -1519 -988 -1503 988
rect -1569 -1000 -1503 -988
rect -1473 988 -1407 1000
rect -1473 -988 -1457 988
rect -1423 -988 -1407 988
rect -1473 -1000 -1407 -988
rect -1377 988 -1311 1000
rect -1377 -988 -1361 988
rect -1327 -988 -1311 988
rect -1377 -1000 -1311 -988
rect -1281 988 -1215 1000
rect -1281 -988 -1265 988
rect -1231 -988 -1215 988
rect -1281 -1000 -1215 -988
rect -1185 988 -1119 1000
rect -1185 -988 -1169 988
rect -1135 -988 -1119 988
rect -1185 -1000 -1119 -988
rect -1089 988 -1023 1000
rect -1089 -988 -1073 988
rect -1039 -988 -1023 988
rect -1089 -1000 -1023 -988
rect -993 988 -927 1000
rect -993 -988 -977 988
rect -943 -988 -927 988
rect -993 -1000 -927 -988
rect -897 988 -831 1000
rect -897 -988 -881 988
rect -847 -988 -831 988
rect -897 -1000 -831 -988
rect -801 988 -735 1000
rect -801 -988 -785 988
rect -751 -988 -735 988
rect -801 -1000 -735 -988
rect -705 988 -639 1000
rect -705 -988 -689 988
rect -655 -988 -639 988
rect -705 -1000 -639 -988
rect -609 988 -543 1000
rect -609 -988 -593 988
rect -559 -988 -543 988
rect -609 -1000 -543 -988
rect -513 988 -447 1000
rect -513 -988 -497 988
rect -463 -988 -447 988
rect -513 -1000 -447 -988
rect -417 988 -351 1000
rect -417 -988 -401 988
rect -367 -988 -351 988
rect -417 -1000 -351 -988
rect -321 988 -255 1000
rect -321 -988 -305 988
rect -271 -988 -255 988
rect -321 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 321 1000
rect 255 -988 271 988
rect 305 -988 321 988
rect 255 -1000 321 -988
rect 351 988 417 1000
rect 351 -988 367 988
rect 401 -988 417 988
rect 351 -1000 417 -988
rect 447 988 513 1000
rect 447 -988 463 988
rect 497 -988 513 988
rect 447 -1000 513 -988
rect 543 988 609 1000
rect 543 -988 559 988
rect 593 -988 609 988
rect 543 -1000 609 -988
rect 639 988 705 1000
rect 639 -988 655 988
rect 689 -988 705 988
rect 639 -1000 705 -988
rect 735 988 801 1000
rect 735 -988 751 988
rect 785 -988 801 988
rect 735 -1000 801 -988
rect 831 988 897 1000
rect 831 -988 847 988
rect 881 -988 897 988
rect 831 -1000 897 -988
rect 927 988 993 1000
rect 927 -988 943 988
rect 977 -988 993 988
rect 927 -1000 993 -988
rect 1023 988 1089 1000
rect 1023 -988 1039 988
rect 1073 -988 1089 988
rect 1023 -1000 1089 -988
rect 1119 988 1185 1000
rect 1119 -988 1135 988
rect 1169 -988 1185 988
rect 1119 -1000 1185 -988
rect 1215 988 1281 1000
rect 1215 -988 1231 988
rect 1265 -988 1281 988
rect 1215 -1000 1281 -988
rect 1311 988 1377 1000
rect 1311 -988 1327 988
rect 1361 -988 1377 988
rect 1311 -1000 1377 -988
rect 1407 988 1473 1000
rect 1407 -988 1423 988
rect 1457 -988 1473 988
rect 1407 -1000 1473 -988
rect 1503 988 1569 1000
rect 1503 -988 1519 988
rect 1553 -988 1569 988
rect 1503 -1000 1569 -988
rect 1599 988 1665 1000
rect 1599 -988 1615 988
rect 1649 -988 1665 988
rect 1599 -1000 1665 -988
rect 1695 988 1761 1000
rect 1695 -988 1711 988
rect 1745 -988 1761 988
rect 1695 -1000 1761 -988
rect 1791 988 1857 1000
rect 1791 -988 1807 988
rect 1841 -988 1857 988
rect 1791 -1000 1857 -988
rect 1887 988 1953 1000
rect 1887 -988 1903 988
rect 1937 -988 1953 988
rect 1887 -1000 1953 -988
rect 1983 988 2049 1000
rect 1983 -988 1999 988
rect 2033 -988 2049 988
rect 1983 -1000 2049 -988
rect 2079 988 2145 1000
rect 2079 -988 2095 988
rect 2129 -988 2145 988
rect 2079 -1000 2145 -988
rect 2175 988 2241 1000
rect 2175 -988 2191 988
rect 2225 -988 2241 988
rect 2175 -1000 2241 -988
rect 2271 988 2337 1000
rect 2271 -988 2287 988
rect 2321 -988 2337 988
rect 2271 -1000 2337 -988
rect 2367 988 2433 1000
rect 2367 -988 2383 988
rect 2417 -988 2433 988
rect 2367 -1000 2433 -988
rect 2463 988 2529 1000
rect 2463 -988 2479 988
rect 2513 -988 2529 988
rect 2463 -1000 2529 -988
rect 2559 988 2625 1000
rect 2559 -988 2575 988
rect 2609 -988 2625 988
rect 2559 -1000 2625 -988
rect 2655 988 2721 1000
rect 2655 -988 2671 988
rect 2705 -988 2721 988
rect 2655 -1000 2721 -988
rect 2751 988 2817 1000
rect 2751 -988 2767 988
rect 2801 -988 2817 988
rect 2751 -1000 2817 -988
rect 2847 988 2909 1000
rect 2847 -988 2863 988
rect 2897 -988 2909 988
rect 2847 -1000 2909 -988
<< ndiffc >>
rect -2897 -988 -2863 988
rect -2801 -988 -2767 988
rect -2705 -988 -2671 988
rect -2609 -988 -2575 988
rect -2513 -988 -2479 988
rect -2417 -988 -2383 988
rect -2321 -988 -2287 988
rect -2225 -988 -2191 988
rect -2129 -988 -2095 988
rect -2033 -988 -1999 988
rect -1937 -988 -1903 988
rect -1841 -988 -1807 988
rect -1745 -988 -1711 988
rect -1649 -988 -1615 988
rect -1553 -988 -1519 988
rect -1457 -988 -1423 988
rect -1361 -988 -1327 988
rect -1265 -988 -1231 988
rect -1169 -988 -1135 988
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
rect 1135 -988 1169 988
rect 1231 -988 1265 988
rect 1327 -988 1361 988
rect 1423 -988 1457 988
rect 1519 -988 1553 988
rect 1615 -988 1649 988
rect 1711 -988 1745 988
rect 1807 -988 1841 988
rect 1903 -988 1937 988
rect 1999 -988 2033 988
rect 2095 -988 2129 988
rect 2191 -988 2225 988
rect 2287 -988 2321 988
rect 2383 -988 2417 988
rect 2479 -988 2513 988
rect 2575 -988 2609 988
rect 2671 -988 2705 988
rect 2767 -988 2801 988
rect 2863 -988 2897 988
<< poly >>
rect -2847 1000 -2817 1026
rect -2751 1000 -2721 1026
rect -2655 1000 -2625 1026
rect -2559 1000 -2529 1026
rect -2463 1000 -2433 1026
rect -2367 1000 -2337 1026
rect -2271 1000 -2241 1026
rect -2175 1000 -2145 1026
rect -2079 1000 -2049 1026
rect -1983 1000 -1953 1026
rect -1887 1000 -1857 1026
rect -1791 1000 -1761 1026
rect -1695 1000 -1665 1026
rect -1599 1000 -1569 1026
rect -1503 1000 -1473 1026
rect -1407 1000 -1377 1026
rect -1311 1000 -1281 1026
rect -1215 1000 -1185 1026
rect -1119 1000 -1089 1026
rect -1023 1000 -993 1026
rect -927 1000 -897 1026
rect -831 1000 -801 1026
rect -735 1000 -705 1026
rect -639 1000 -609 1026
rect -543 1000 -513 1026
rect -447 1000 -417 1026
rect -351 1000 -321 1026
rect -255 1000 -225 1026
rect -159 1000 -129 1026
rect -63 1000 -33 1026
rect 33 1000 63 1026
rect 129 1000 159 1026
rect 225 1000 255 1026
rect 321 1000 351 1026
rect 417 1000 447 1026
rect 513 1000 543 1026
rect 609 1000 639 1026
rect 705 1000 735 1026
rect 801 1000 831 1026
rect 897 1000 927 1026
rect 993 1000 1023 1026
rect 1089 1000 1119 1026
rect 1185 1000 1215 1026
rect 1281 1000 1311 1026
rect 1377 1000 1407 1026
rect 1473 1000 1503 1026
rect 1569 1000 1599 1026
rect 1665 1000 1695 1026
rect 1761 1000 1791 1026
rect 1857 1000 1887 1026
rect 1953 1000 1983 1026
rect 2049 1000 2079 1026
rect 2145 1000 2175 1026
rect 2241 1000 2271 1026
rect 2337 1000 2367 1026
rect 2433 1000 2463 1026
rect 2529 1000 2559 1026
rect 2625 1000 2655 1026
rect 2721 1000 2751 1026
rect 2817 1000 2847 1026
rect -2847 -1020 -2817 -1000
rect -2751 -1020 -2721 -1000
rect -2655 -1020 -2625 -1000
rect -2559 -1020 -2529 -1000
rect -2463 -1020 -2433 -1000
rect -2367 -1020 -2337 -1000
rect -2271 -1020 -2241 -1000
rect -2175 -1020 -2145 -1000
rect -2079 -1020 -2049 -1000
rect -1983 -1020 -1953 -1000
rect -1887 -1020 -1857 -1000
rect -1791 -1020 -1761 -1000
rect -1695 -1020 -1665 -1000
rect -1599 -1020 -1569 -1000
rect -1503 -1020 -1473 -1000
rect -1407 -1020 -1377 -1000
rect -1311 -1020 -1281 -1000
rect -1215 -1020 -1185 -1000
rect -1119 -1020 -1089 -1000
rect -1023 -1020 -993 -1000
rect -927 -1020 -897 -1000
rect -831 -1020 -801 -1000
rect -735 -1020 -705 -1000
rect -639 -1020 -609 -1000
rect -543 -1020 -513 -1000
rect -447 -1020 -417 -1000
rect -351 -1020 -321 -1000
rect -255 -1020 -225 -1000
rect -159 -1020 -129 -1000
rect -63 -1020 -33 -1000
rect 33 -1020 63 -1000
rect 129 -1020 159 -1000
rect 225 -1020 255 -1000
rect 321 -1020 351 -1000
rect 417 -1020 447 -1000
rect 513 -1020 543 -1000
rect 609 -1020 639 -1000
rect 705 -1020 735 -1000
rect 801 -1020 831 -1000
rect 897 -1020 927 -1000
rect 993 -1020 1023 -1000
rect 1089 -1020 1119 -1000
rect 1185 -1020 1215 -1000
rect 1281 -1020 1311 -1000
rect 1377 -1020 1407 -1000
rect 1473 -1020 1503 -1000
rect 1569 -1020 1599 -1000
rect 1665 -1020 1695 -1000
rect 1761 -1020 1791 -1000
rect 1857 -1020 1887 -1000
rect 1953 -1020 1983 -1000
rect 2049 -1020 2079 -1000
rect 2145 -1020 2175 -1000
rect 2241 -1020 2271 -1000
rect 2337 -1020 2367 -1000
rect 2433 -1020 2463 -1000
rect 2529 -1020 2559 -1000
rect 2625 -1020 2655 -1000
rect 2721 -1020 2751 -1000
rect 2817 -1020 2847 -1000
rect -2883 -1038 2909 -1020
rect -2883 -1072 -2849 -1038
rect -2815 -1072 -2657 -1038
rect -2623 -1072 -2465 -1038
rect -2431 -1072 -2273 -1038
rect -2239 -1072 -2081 -1038
rect -2047 -1072 -1889 -1038
rect -1855 -1072 -1697 -1038
rect -1663 -1072 -1505 -1038
rect -1471 -1072 -1313 -1038
rect -1279 -1072 -1121 -1038
rect -1087 -1072 -929 -1038
rect -895 -1072 -737 -1038
rect -703 -1072 -545 -1038
rect -511 -1072 -353 -1038
rect -319 -1072 -161 -1038
rect -127 -1072 31 -1038
rect 65 -1072 223 -1038
rect 257 -1072 415 -1038
rect 449 -1072 607 -1038
rect 641 -1072 799 -1038
rect 833 -1072 991 -1038
rect 1025 -1072 1183 -1038
rect 1217 -1072 1375 -1038
rect 1409 -1072 1567 -1038
rect 1601 -1072 1759 -1038
rect 1793 -1072 1951 -1038
rect 1985 -1072 2143 -1038
rect 2177 -1072 2335 -1038
rect 2369 -1072 2527 -1038
rect 2561 -1072 2719 -1038
rect 2753 -1072 2909 -1038
rect -2883 -1088 2909 -1072
<< polycont >>
rect -2849 -1072 -2815 -1038
rect -2657 -1072 -2623 -1038
rect -2465 -1072 -2431 -1038
rect -2273 -1072 -2239 -1038
rect -2081 -1072 -2047 -1038
rect -1889 -1072 -1855 -1038
rect -1697 -1072 -1663 -1038
rect -1505 -1072 -1471 -1038
rect -1313 -1072 -1279 -1038
rect -1121 -1072 -1087 -1038
rect -929 -1072 -895 -1038
rect -737 -1072 -703 -1038
rect -545 -1072 -511 -1038
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
rect 415 -1072 449 -1038
rect 607 -1072 641 -1038
rect 799 -1072 833 -1038
rect 991 -1072 1025 -1038
rect 1183 -1072 1217 -1038
rect 1375 -1072 1409 -1038
rect 1567 -1072 1601 -1038
rect 1759 -1072 1793 -1038
rect 1951 -1072 1985 -1038
rect 2143 -1072 2177 -1038
rect 2335 -1072 2369 -1038
rect 2527 -1072 2561 -1038
rect 2719 -1072 2753 -1038
<< locali >>
rect -2897 988 -2863 1004
rect -2897 -1004 -2863 -988
rect -2801 988 -2767 1004
rect -2801 -1004 -2767 -988
rect -2705 988 -2671 1004
rect -2705 -1004 -2671 -988
rect -2609 988 -2575 1004
rect -2609 -1004 -2575 -988
rect -2513 988 -2479 1004
rect -2513 -1004 -2479 -988
rect -2417 988 -2383 1004
rect -2417 -1004 -2383 -988
rect -2321 988 -2287 1004
rect -2321 -1004 -2287 -988
rect -2225 988 -2191 1004
rect -2225 -1004 -2191 -988
rect -2129 988 -2095 1004
rect -2129 -1004 -2095 -988
rect -2033 988 -1999 1004
rect -2033 -1004 -1999 -988
rect -1937 988 -1903 1004
rect -1937 -1004 -1903 -988
rect -1841 988 -1807 1004
rect -1841 -1004 -1807 -988
rect -1745 988 -1711 1004
rect -1745 -1004 -1711 -988
rect -1649 988 -1615 1004
rect -1649 -1004 -1615 -988
rect -1553 988 -1519 1004
rect -1553 -1004 -1519 -988
rect -1457 988 -1423 1004
rect -1457 -1004 -1423 -988
rect -1361 988 -1327 1004
rect -1361 -1004 -1327 -988
rect -1265 988 -1231 1004
rect -1265 -1004 -1231 -988
rect -1169 988 -1135 1004
rect -1169 -1004 -1135 -988
rect -1073 988 -1039 1004
rect -1073 -1004 -1039 -988
rect -977 988 -943 1004
rect -977 -1004 -943 -988
rect -881 988 -847 1004
rect -881 -1004 -847 -988
rect -785 988 -751 1004
rect -785 -1004 -751 -988
rect -689 988 -655 1004
rect -689 -1004 -655 -988
rect -593 988 -559 1004
rect -593 -1004 -559 -988
rect -497 988 -463 1004
rect -497 -1004 -463 -988
rect -401 988 -367 1004
rect -401 -1004 -367 -988
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect 367 988 401 1004
rect 367 -1004 401 -988
rect 463 988 497 1004
rect 463 -1004 497 -988
rect 559 988 593 1004
rect 559 -1004 593 -988
rect 655 988 689 1004
rect 655 -1004 689 -988
rect 751 988 785 1004
rect 751 -1004 785 -988
rect 847 988 881 1004
rect 847 -1004 881 -988
rect 943 988 977 1004
rect 943 -1004 977 -988
rect 1039 988 1073 1004
rect 1039 -1004 1073 -988
rect 1135 988 1169 1004
rect 1135 -1004 1169 -988
rect 1231 988 1265 1004
rect 1231 -1004 1265 -988
rect 1327 988 1361 1004
rect 1327 -1004 1361 -988
rect 1423 988 1457 1004
rect 1423 -1004 1457 -988
rect 1519 988 1553 1004
rect 1519 -1004 1553 -988
rect 1615 988 1649 1004
rect 1615 -1004 1649 -988
rect 1711 988 1745 1004
rect 1711 -1004 1745 -988
rect 1807 988 1841 1004
rect 1807 -1004 1841 -988
rect 1903 988 1937 1004
rect 1903 -1004 1937 -988
rect 1999 988 2033 1004
rect 1999 -1004 2033 -988
rect 2095 988 2129 1004
rect 2095 -1004 2129 -988
rect 2191 988 2225 1004
rect 2191 -1004 2225 -988
rect 2287 988 2321 1004
rect 2287 -1004 2321 -988
rect 2383 988 2417 1004
rect 2383 -1004 2417 -988
rect 2479 988 2513 1004
rect 2479 -1004 2513 -988
rect 2575 988 2609 1004
rect 2575 -1004 2609 -988
rect 2671 988 2705 1004
rect 2671 -1004 2705 -988
rect 2767 988 2801 1004
rect 2767 -1004 2801 -988
rect 2863 988 2897 1004
rect 2863 -1004 2897 -988
rect -2865 -1072 -2849 -1038
rect -2815 -1072 -2799 -1038
rect -2673 -1072 -2657 -1038
rect -2623 -1072 -2607 -1038
rect -2481 -1072 -2465 -1038
rect -2431 -1072 -2415 -1038
rect -2289 -1072 -2273 -1038
rect -2239 -1072 -2223 -1038
rect -2097 -1072 -2081 -1038
rect -2047 -1072 -2031 -1038
rect -1905 -1072 -1889 -1038
rect -1855 -1072 -1839 -1038
rect -1713 -1072 -1697 -1038
rect -1663 -1072 -1647 -1038
rect -1521 -1072 -1505 -1038
rect -1471 -1072 -1455 -1038
rect -1329 -1072 -1313 -1038
rect -1279 -1072 -1263 -1038
rect -1137 -1072 -1121 -1038
rect -1087 -1072 -1071 -1038
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect 975 -1072 991 -1038
rect 1025 -1072 1041 -1038
rect 1167 -1072 1183 -1038
rect 1217 -1072 1233 -1038
rect 1359 -1072 1375 -1038
rect 1409 -1072 1425 -1038
rect 1551 -1072 1567 -1038
rect 1601 -1072 1617 -1038
rect 1743 -1072 1759 -1038
rect 1793 -1072 1809 -1038
rect 1935 -1072 1951 -1038
rect 1985 -1072 2001 -1038
rect 2127 -1072 2143 -1038
rect 2177 -1072 2193 -1038
rect 2319 -1072 2335 -1038
rect 2369 -1072 2385 -1038
rect 2511 -1072 2527 -1038
rect 2561 -1072 2577 -1038
rect 2703 -1072 2719 -1038
rect 2753 -1072 2769 -1038
<< viali >>
rect -2897 -988 -2863 988
rect -2801 -988 -2767 988
rect -2705 -988 -2671 988
rect -2609 -988 -2575 988
rect -2513 -988 -2479 988
rect -2417 -988 -2383 988
rect -2321 -988 -2287 988
rect -2225 -988 -2191 988
rect -2129 -988 -2095 988
rect -2033 -988 -1999 988
rect -1937 -988 -1903 988
rect -1841 -988 -1807 988
rect -1745 -988 -1711 988
rect -1649 -988 -1615 988
rect -1553 -988 -1519 988
rect -1457 -988 -1423 988
rect -1361 -988 -1327 988
rect -1265 -988 -1231 988
rect -1169 -988 -1135 988
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
rect 1135 -988 1169 988
rect 1231 -988 1265 988
rect 1327 -988 1361 988
rect 1423 -988 1457 988
rect 1519 -988 1553 988
rect 1615 -988 1649 988
rect 1711 -988 1745 988
rect 1807 -988 1841 988
rect 1903 -988 1937 988
rect 1999 -988 2033 988
rect 2095 -988 2129 988
rect 2191 -988 2225 988
rect 2287 -988 2321 988
rect 2383 -988 2417 988
rect 2479 -988 2513 988
rect 2575 -988 2609 988
rect 2671 -988 2705 988
rect 2767 -988 2801 988
rect 2863 -988 2897 988
rect -2849 -1072 -2815 -1038
rect -2657 -1072 -2623 -1038
rect -2465 -1072 -2431 -1038
rect -2273 -1072 -2239 -1038
rect -2081 -1072 -2047 -1038
rect -1889 -1072 -1855 -1038
rect -1697 -1072 -1663 -1038
rect -1505 -1072 -1471 -1038
rect -1313 -1072 -1279 -1038
rect -1121 -1072 -1087 -1038
rect -929 -1072 -895 -1038
rect -737 -1072 -703 -1038
rect -545 -1072 -511 -1038
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
rect 415 -1072 449 -1038
rect 607 -1072 641 -1038
rect 799 -1072 833 -1038
rect 991 -1072 1025 -1038
rect 1183 -1072 1217 -1038
rect 1375 -1072 1409 -1038
rect 1567 -1072 1601 -1038
rect 1759 -1072 1793 -1038
rect 1951 -1072 1985 -1038
rect 2143 -1072 2177 -1038
rect 2335 -1072 2369 -1038
rect 2527 -1072 2561 -1038
rect 2719 -1072 2753 -1038
<< metal1 >>
rect -2903 988 -2857 1000
rect -2903 -988 -2897 988
rect -2863 -988 -2857 988
rect -2903 -1000 -2857 -988
rect -2807 988 -2761 1000
rect -2807 -988 -2801 988
rect -2767 -988 -2761 988
rect -2807 -1000 -2761 -988
rect -2711 988 -2665 1000
rect -2711 -988 -2705 988
rect -2671 -988 -2665 988
rect -2711 -1000 -2665 -988
rect -2615 988 -2569 1000
rect -2615 -988 -2609 988
rect -2575 -988 -2569 988
rect -2615 -1000 -2569 -988
rect -2519 988 -2473 1000
rect -2519 -988 -2513 988
rect -2479 -988 -2473 988
rect -2519 -1000 -2473 -988
rect -2423 988 -2377 1000
rect -2423 -988 -2417 988
rect -2383 -988 -2377 988
rect -2423 -1000 -2377 -988
rect -2327 988 -2281 1000
rect -2327 -988 -2321 988
rect -2287 -988 -2281 988
rect -2327 -1000 -2281 -988
rect -2231 988 -2185 1000
rect -2231 -988 -2225 988
rect -2191 -988 -2185 988
rect -2231 -1000 -2185 -988
rect -2135 988 -2089 1000
rect -2135 -988 -2129 988
rect -2095 -988 -2089 988
rect -2135 -1000 -2089 -988
rect -2039 988 -1993 1000
rect -2039 -988 -2033 988
rect -1999 -988 -1993 988
rect -2039 -1000 -1993 -988
rect -1943 988 -1897 1000
rect -1943 -988 -1937 988
rect -1903 -988 -1897 988
rect -1943 -1000 -1897 -988
rect -1847 988 -1801 1000
rect -1847 -988 -1841 988
rect -1807 -988 -1801 988
rect -1847 -1000 -1801 -988
rect -1751 988 -1705 1000
rect -1751 -988 -1745 988
rect -1711 -988 -1705 988
rect -1751 -1000 -1705 -988
rect -1655 988 -1609 1000
rect -1655 -988 -1649 988
rect -1615 -988 -1609 988
rect -1655 -1000 -1609 -988
rect -1559 988 -1513 1000
rect -1559 -988 -1553 988
rect -1519 -988 -1513 988
rect -1559 -1000 -1513 -988
rect -1463 988 -1417 1000
rect -1463 -988 -1457 988
rect -1423 -988 -1417 988
rect -1463 -1000 -1417 -988
rect -1367 988 -1321 1000
rect -1367 -988 -1361 988
rect -1327 -988 -1321 988
rect -1367 -1000 -1321 -988
rect -1271 988 -1225 1000
rect -1271 -988 -1265 988
rect -1231 -988 -1225 988
rect -1271 -1000 -1225 -988
rect -1175 988 -1129 1000
rect -1175 -988 -1169 988
rect -1135 -988 -1129 988
rect -1175 -1000 -1129 -988
rect -1079 988 -1033 1000
rect -1079 -988 -1073 988
rect -1039 -988 -1033 988
rect -1079 -1000 -1033 -988
rect -983 988 -937 1000
rect -983 -988 -977 988
rect -943 -988 -937 988
rect -983 -1000 -937 -988
rect -887 988 -841 1000
rect -887 -988 -881 988
rect -847 -988 -841 988
rect -887 -1000 -841 -988
rect -791 988 -745 1000
rect -791 -988 -785 988
rect -751 -988 -745 988
rect -791 -1000 -745 -988
rect -695 988 -649 1000
rect -695 -988 -689 988
rect -655 -988 -649 988
rect -695 -1000 -649 -988
rect -599 988 -553 1000
rect -599 -988 -593 988
rect -559 -988 -553 988
rect -599 -1000 -553 -988
rect -503 988 -457 1000
rect -503 -988 -497 988
rect -463 -988 -457 988
rect -503 -1000 -457 -988
rect -407 988 -361 1000
rect -407 -988 -401 988
rect -367 -988 -361 988
rect -407 -1000 -361 -988
rect -311 988 -265 1000
rect -311 -988 -305 988
rect -271 -988 -265 988
rect -311 -1000 -265 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 265 988 311 1000
rect 265 -988 271 988
rect 305 -988 311 988
rect 265 -1000 311 -988
rect 361 988 407 1000
rect 361 -988 367 988
rect 401 -988 407 988
rect 361 -1000 407 -988
rect 457 988 503 1000
rect 457 -988 463 988
rect 497 -988 503 988
rect 457 -1000 503 -988
rect 553 988 599 1000
rect 553 -988 559 988
rect 593 -988 599 988
rect 553 -1000 599 -988
rect 649 988 695 1000
rect 649 -988 655 988
rect 689 -988 695 988
rect 649 -1000 695 -988
rect 745 988 791 1000
rect 745 -988 751 988
rect 785 -988 791 988
rect 745 -1000 791 -988
rect 841 988 887 1000
rect 841 -988 847 988
rect 881 -988 887 988
rect 841 -1000 887 -988
rect 937 988 983 1000
rect 937 -988 943 988
rect 977 -988 983 988
rect 937 -1000 983 -988
rect 1033 988 1079 1000
rect 1033 -988 1039 988
rect 1073 -988 1079 988
rect 1033 -1000 1079 -988
rect 1129 988 1175 1000
rect 1129 -988 1135 988
rect 1169 -988 1175 988
rect 1129 -1000 1175 -988
rect 1225 988 1271 1000
rect 1225 -988 1231 988
rect 1265 -988 1271 988
rect 1225 -1000 1271 -988
rect 1321 988 1367 1000
rect 1321 -988 1327 988
rect 1361 -988 1367 988
rect 1321 -1000 1367 -988
rect 1417 988 1463 1000
rect 1417 -988 1423 988
rect 1457 -988 1463 988
rect 1417 -1000 1463 -988
rect 1513 988 1559 1000
rect 1513 -988 1519 988
rect 1553 -988 1559 988
rect 1513 -1000 1559 -988
rect 1609 988 1655 1000
rect 1609 -988 1615 988
rect 1649 -988 1655 988
rect 1609 -1000 1655 -988
rect 1705 988 1751 1000
rect 1705 -988 1711 988
rect 1745 -988 1751 988
rect 1705 -1000 1751 -988
rect 1801 988 1847 1000
rect 1801 -988 1807 988
rect 1841 -988 1847 988
rect 1801 -1000 1847 -988
rect 1897 988 1943 1000
rect 1897 -988 1903 988
rect 1937 -988 1943 988
rect 1897 -1000 1943 -988
rect 1993 988 2039 1000
rect 1993 -988 1999 988
rect 2033 -988 2039 988
rect 1993 -1000 2039 -988
rect 2089 988 2135 1000
rect 2089 -988 2095 988
rect 2129 -988 2135 988
rect 2089 -1000 2135 -988
rect 2185 988 2231 1000
rect 2185 -988 2191 988
rect 2225 -988 2231 988
rect 2185 -1000 2231 -988
rect 2281 988 2327 1000
rect 2281 -988 2287 988
rect 2321 -988 2327 988
rect 2281 -1000 2327 -988
rect 2377 988 2423 1000
rect 2377 -988 2383 988
rect 2417 -988 2423 988
rect 2377 -1000 2423 -988
rect 2473 988 2519 1000
rect 2473 -988 2479 988
rect 2513 -988 2519 988
rect 2473 -1000 2519 -988
rect 2569 988 2615 1000
rect 2569 -988 2575 988
rect 2609 -988 2615 988
rect 2569 -1000 2615 -988
rect 2665 988 2711 1000
rect 2665 -988 2671 988
rect 2705 -988 2711 988
rect 2665 -1000 2711 -988
rect 2761 988 2807 1000
rect 2761 -988 2767 988
rect 2801 -988 2807 988
rect 2761 -1000 2807 -988
rect 2857 988 2903 1000
rect 2857 -988 2863 988
rect 2897 -988 2903 988
rect 2857 -1000 2903 -988
rect -2883 -1038 2797 -1030
rect -2883 -1072 -2849 -1038
rect -2815 -1072 -2657 -1038
rect -2623 -1072 -2465 -1038
rect -2431 -1072 -2273 -1038
rect -2239 -1072 -2081 -1038
rect -2047 -1072 -1889 -1038
rect -1855 -1072 -1697 -1038
rect -1663 -1072 -1505 -1038
rect -1471 -1072 -1313 -1038
rect -1279 -1072 -1121 -1038
rect -1087 -1072 -929 -1038
rect -895 -1072 -737 -1038
rect -703 -1072 -545 -1038
rect -511 -1072 -353 -1038
rect -319 -1072 -161 -1038
rect -127 -1072 31 -1038
rect 65 -1072 223 -1038
rect 257 -1072 415 -1038
rect 449 -1072 607 -1038
rect 641 -1072 799 -1038
rect 833 -1072 991 -1038
rect 1025 -1072 1183 -1038
rect 1217 -1072 1375 -1038
rect 1409 -1072 1567 -1038
rect 1601 -1072 1759 -1038
rect 1793 -1072 1951 -1038
rect 1985 -1072 2143 -1038
rect 2177 -1072 2335 -1038
rect 2369 -1072 2527 -1038
rect 2561 -1072 2719 -1038
rect 2753 -1072 2797 -1038
rect -2883 -1088 2797 -1072
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.150 m 1 nf 60 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
