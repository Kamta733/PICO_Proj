** sch_path: /foss/designs/untitled.sch
**.subckt untitled CKS VP VN
*.ipin CKS
*.ipin VP
*.ipin VN
XM1 VP CKS VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=60 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.end
