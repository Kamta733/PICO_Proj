* NGSPICE file created from NmosF29.ext - technology: sky130A

.subckt NmosF29
X0 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=1.048e+14p pd=6.5048e+08u as=9.9e+13p ps=6.099e+08u w=2e+07u l=150000u
X1 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=1.98e+14p pd=1.2198e+09u as=2.038e+14p ps=1.26038e+09u w=2e+07u l=150000u
X2 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X3 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X4 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X5 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X6 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X7 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X8 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X9 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X10 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X11 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X12 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X13 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X14 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X15 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X16 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X17 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X18 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X19 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X20 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X21 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X22 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X23 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X24 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X25 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X26 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X27 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X28 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X29 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X30 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X31 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X32 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X33 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X34 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X35 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X36 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X37 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X38 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X39 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X40 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X41 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X42 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X43 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X44 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X45 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X46 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X47 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X48 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X49 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X50 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X51 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X52 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X53 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X54 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X55 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X56 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X57 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X58 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X59 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X60 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X61 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X62 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X63 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X64 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X65 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X66 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X67 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X68 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X69 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X70 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X71 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X72 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X73 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X74 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X75 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X76 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X77 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X78 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X79 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X80 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X81 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X82 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X83 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X84 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X85 VX OUT OUT OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X86 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X87 VX CKS VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X88 VN CKS VX VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X89 OUT OUT VX OUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
.ends

