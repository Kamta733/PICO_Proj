magic
tech sky130A
timestamp 1661682518
<< nmos >>
rect -35 150 -20 1150
rect 9 150 24 1150
rect 54 150 69 1150
rect 99 150 114 1150
rect 144 150 159 1150
rect 189 150 204 1150
rect 234 150 249 1150
rect 279 150 294 1150
rect 325 150 340 1150
rect 369 150 384 1150
rect 414 150 429 1150
rect 459 150 474 1150
rect 504 150 519 1150
rect 549 150 564 1150
rect 594 150 609 1150
rect 639 150 654 1150
rect 684 150 699 1150
rect 728 150 743 1150
rect 773 150 788 1150
rect 818 150 833 1150
rect 863 150 878 1150
rect 908 150 923 1150
rect 953 150 968 1150
rect 998 150 1013 1150
rect 1044 150 1059 1150
rect 1088 150 1103 1150
rect 1133 150 1148 1150
rect 1178 150 1193 1150
rect 1223 150 1238 1150
rect 1268 150 1283 1150
rect 1313 150 1328 1150
rect 1358 150 1373 1150
rect 1403 150 1418 1150
rect 1447 150 1462 1150
rect 1492 150 1507 1150
rect 1537 150 1552 1150
rect 1582 150 1597 1150
rect 1627 150 1642 1150
rect 1672 150 1687 1150
rect 1717 150 1732 1150
rect 1763 150 1778 1150
rect 1807 150 1822 1150
rect 1852 150 1867 1150
rect 1897 150 1912 1150
rect 1942 150 1957 1150
rect 1987 150 2002 1150
rect 2032 150 2047 1150
rect 2077 150 2092 1150
rect 2122 150 2137 1150
rect 2166 150 2181 1150
rect 2211 150 2226 1150
rect 2256 150 2271 1150
rect 2301 150 2316 1150
rect 2346 150 2361 1150
rect 2391 150 2406 1150
rect 2436 150 2451 1150
rect 2482 150 2497 1150
rect 2526 150 2541 1150
rect 2571 150 2586 1150
rect 2616 150 2631 1150
<< ndiff >>
rect -64 1135 -35 1150
rect -64 1118 -59 1135
rect -42 1118 -35 1135
rect -64 1101 -35 1118
rect -64 1084 -59 1101
rect -42 1084 -35 1101
rect -64 1067 -35 1084
rect -64 1050 -59 1067
rect -42 1050 -35 1067
rect -64 1033 -35 1050
rect -64 1016 -59 1033
rect -42 1016 -35 1033
rect -64 999 -35 1016
rect -64 982 -58 999
rect -41 982 -35 999
rect -64 965 -35 982
rect -64 948 -58 965
rect -41 948 -35 965
rect -64 931 -35 948
rect -64 914 -58 931
rect -41 914 -35 931
rect -64 897 -35 914
rect -64 880 -58 897
rect -41 880 -35 897
rect -64 863 -35 880
rect -64 846 -58 863
rect -41 846 -35 863
rect -64 829 -35 846
rect -64 812 -58 829
rect -41 812 -35 829
rect -64 795 -35 812
rect -64 778 -58 795
rect -41 778 -35 795
rect -64 761 -35 778
rect -64 744 -58 761
rect -41 744 -35 761
rect -64 727 -35 744
rect -64 710 -58 727
rect -41 710 -35 727
rect -64 693 -35 710
rect -64 676 -58 693
rect -41 676 -35 693
rect -64 659 -35 676
rect -64 642 -58 659
rect -41 642 -35 659
rect -64 625 -35 642
rect -64 608 -58 625
rect -41 608 -35 625
rect -64 591 -35 608
rect -64 574 -58 591
rect -41 574 -35 591
rect -64 557 -35 574
rect -64 540 -58 557
rect -41 540 -35 557
rect -64 523 -35 540
rect -64 506 -58 523
rect -41 506 -35 523
rect -64 489 -35 506
rect -64 472 -58 489
rect -41 472 -35 489
rect -64 455 -35 472
rect -64 438 -58 455
rect -41 438 -35 455
rect -64 421 -35 438
rect -64 404 -58 421
rect -41 404 -35 421
rect -64 387 -35 404
rect -64 370 -58 387
rect -41 370 -35 387
rect -64 353 -35 370
rect -64 336 -58 353
rect -41 336 -35 353
rect -64 319 -35 336
rect -64 302 -58 319
rect -41 302 -35 319
rect -64 285 -35 302
rect -64 268 -58 285
rect -41 268 -35 285
rect -64 251 -35 268
rect -64 234 -58 251
rect -41 234 -35 251
rect -64 217 -35 234
rect -64 200 -58 217
rect -41 200 -35 217
rect -64 183 -35 200
rect -64 166 -58 183
rect -41 166 -35 183
rect -64 150 -35 166
rect -20 1137 9 1150
rect -20 1120 -14 1137
rect 3 1120 9 1137
rect -20 1103 9 1120
rect -20 1086 -14 1103
rect 3 1086 9 1103
rect -20 1069 9 1086
rect -20 1052 -14 1069
rect 3 1052 9 1069
rect -20 1035 9 1052
rect -20 1018 -14 1035
rect 3 1018 9 1035
rect -20 1001 9 1018
rect -20 984 -14 1001
rect 3 984 9 1001
rect -20 967 9 984
rect -20 950 -14 967
rect 3 950 9 967
rect -20 933 9 950
rect -20 916 -14 933
rect 3 916 9 933
rect -20 899 9 916
rect -20 882 -14 899
rect 3 882 9 899
rect -20 865 9 882
rect -20 848 -14 865
rect 3 848 9 865
rect -20 831 9 848
rect -20 814 -14 831
rect 3 814 9 831
rect -20 797 9 814
rect -20 780 -14 797
rect 3 780 9 797
rect -20 763 9 780
rect -20 746 -14 763
rect 3 746 9 763
rect -20 729 9 746
rect -20 712 -14 729
rect 3 712 9 729
rect -20 695 9 712
rect -20 678 -14 695
rect 3 678 9 695
rect -20 661 9 678
rect -20 644 -14 661
rect 3 644 9 661
rect -20 627 9 644
rect -20 610 -14 627
rect 3 610 9 627
rect -20 593 9 610
rect -20 576 -14 593
rect 3 576 9 593
rect -20 559 9 576
rect -20 542 -14 559
rect 3 542 9 559
rect -20 525 9 542
rect -20 508 -14 525
rect 3 508 9 525
rect -20 491 9 508
rect -20 474 -14 491
rect 3 474 9 491
rect -20 457 9 474
rect -20 440 -14 457
rect 3 440 9 457
rect -20 423 9 440
rect -20 406 -14 423
rect 3 406 9 423
rect -20 389 9 406
rect -20 372 -14 389
rect 3 372 9 389
rect -20 355 9 372
rect -20 338 -14 355
rect 3 338 9 355
rect -20 321 9 338
rect -20 304 -14 321
rect 3 304 9 321
rect -20 287 9 304
rect -20 270 -14 287
rect 3 270 9 287
rect -20 253 9 270
rect -20 236 -14 253
rect 3 236 9 253
rect -20 219 9 236
rect -20 202 -14 219
rect 3 202 9 219
rect -20 185 9 202
rect -20 168 -14 185
rect 3 168 9 185
rect -20 150 9 168
rect 24 1135 54 1150
rect 24 1118 30 1135
rect 47 1118 54 1135
rect 24 1101 54 1118
rect 24 1084 30 1101
rect 47 1084 54 1101
rect 24 1067 54 1084
rect 24 1050 30 1067
rect 47 1050 54 1067
rect 24 1033 54 1050
rect 24 1016 30 1033
rect 47 1016 54 1033
rect 24 999 54 1016
rect 24 982 31 999
rect 48 982 54 999
rect 24 965 54 982
rect 24 948 31 965
rect 48 948 54 965
rect 24 931 54 948
rect 24 914 31 931
rect 48 914 54 931
rect 24 897 54 914
rect 24 880 31 897
rect 48 880 54 897
rect 24 863 54 880
rect 24 846 31 863
rect 48 846 54 863
rect 24 829 54 846
rect 24 812 31 829
rect 48 812 54 829
rect 24 795 54 812
rect 24 778 31 795
rect 48 778 54 795
rect 24 761 54 778
rect 24 744 31 761
rect 48 744 54 761
rect 24 727 54 744
rect 24 710 31 727
rect 48 710 54 727
rect 24 693 54 710
rect 24 676 31 693
rect 48 676 54 693
rect 24 659 54 676
rect 24 642 31 659
rect 48 642 54 659
rect 24 625 54 642
rect 24 608 31 625
rect 48 608 54 625
rect 24 591 54 608
rect 24 574 31 591
rect 48 574 54 591
rect 24 557 54 574
rect 24 540 31 557
rect 48 540 54 557
rect 24 523 54 540
rect 24 506 31 523
rect 48 506 54 523
rect 24 489 54 506
rect 24 472 31 489
rect 48 472 54 489
rect 24 455 54 472
rect 24 438 31 455
rect 48 438 54 455
rect 24 421 54 438
rect 24 404 31 421
rect 48 404 54 421
rect 24 387 54 404
rect 24 370 31 387
rect 48 370 54 387
rect 24 353 54 370
rect 24 336 31 353
rect 48 336 54 353
rect 24 319 54 336
rect 24 302 31 319
rect 48 302 54 319
rect 24 285 54 302
rect 24 268 31 285
rect 48 268 54 285
rect 24 251 54 268
rect 24 234 31 251
rect 48 234 54 251
rect 24 217 54 234
rect 24 200 31 217
rect 48 200 54 217
rect 24 183 54 200
rect 24 166 31 183
rect 48 166 54 183
rect 24 150 54 166
rect 69 1135 99 1150
rect 69 1118 75 1135
rect 92 1118 99 1135
rect 69 1101 99 1118
rect 69 1084 75 1101
rect 92 1084 99 1101
rect 69 1067 99 1084
rect 69 1050 75 1067
rect 92 1050 99 1067
rect 69 1033 99 1050
rect 69 1016 75 1033
rect 92 1016 99 1033
rect 69 999 99 1016
rect 69 982 76 999
rect 93 982 99 999
rect 69 965 99 982
rect 69 948 76 965
rect 93 948 99 965
rect 69 931 99 948
rect 69 914 76 931
rect 93 914 99 931
rect 69 897 99 914
rect 69 880 76 897
rect 93 880 99 897
rect 69 863 99 880
rect 69 846 76 863
rect 93 846 99 863
rect 69 829 99 846
rect 69 812 76 829
rect 93 812 99 829
rect 69 795 99 812
rect 69 778 76 795
rect 93 778 99 795
rect 69 761 99 778
rect 69 744 76 761
rect 93 744 99 761
rect 69 727 99 744
rect 69 710 76 727
rect 93 710 99 727
rect 69 693 99 710
rect 69 676 76 693
rect 93 676 99 693
rect 69 659 99 676
rect 69 642 76 659
rect 93 642 99 659
rect 69 625 99 642
rect 69 608 76 625
rect 93 608 99 625
rect 69 591 99 608
rect 69 574 76 591
rect 93 574 99 591
rect 69 557 99 574
rect 69 540 76 557
rect 93 540 99 557
rect 69 523 99 540
rect 69 506 76 523
rect 93 506 99 523
rect 69 489 99 506
rect 69 472 76 489
rect 93 472 99 489
rect 69 455 99 472
rect 69 438 76 455
rect 93 438 99 455
rect 69 421 99 438
rect 69 404 76 421
rect 93 404 99 421
rect 69 387 99 404
rect 69 370 76 387
rect 93 370 99 387
rect 69 353 99 370
rect 69 336 76 353
rect 93 336 99 353
rect 69 319 99 336
rect 69 302 76 319
rect 93 302 99 319
rect 69 285 99 302
rect 69 268 76 285
rect 93 268 99 285
rect 69 251 99 268
rect 69 234 76 251
rect 93 234 99 251
rect 69 217 99 234
rect 69 200 76 217
rect 93 200 99 217
rect 69 183 99 200
rect 69 166 76 183
rect 93 166 99 183
rect 69 150 99 166
rect 114 1135 144 1150
rect 114 1118 120 1135
rect 137 1118 144 1135
rect 114 1101 144 1118
rect 114 1084 120 1101
rect 137 1084 144 1101
rect 114 1067 144 1084
rect 114 1050 120 1067
rect 137 1050 144 1067
rect 114 1033 144 1050
rect 114 1016 120 1033
rect 137 1016 144 1033
rect 114 999 144 1016
rect 114 982 121 999
rect 138 982 144 999
rect 114 965 144 982
rect 114 948 121 965
rect 138 948 144 965
rect 114 931 144 948
rect 114 914 121 931
rect 138 914 144 931
rect 114 897 144 914
rect 114 880 121 897
rect 138 880 144 897
rect 114 863 144 880
rect 114 846 121 863
rect 138 846 144 863
rect 114 829 144 846
rect 114 812 121 829
rect 138 812 144 829
rect 114 795 144 812
rect 114 778 121 795
rect 138 778 144 795
rect 114 761 144 778
rect 114 744 121 761
rect 138 744 144 761
rect 114 727 144 744
rect 114 710 121 727
rect 138 710 144 727
rect 114 693 144 710
rect 114 676 121 693
rect 138 676 144 693
rect 114 659 144 676
rect 114 642 121 659
rect 138 642 144 659
rect 114 625 144 642
rect 114 608 121 625
rect 138 608 144 625
rect 114 591 144 608
rect 114 574 121 591
rect 138 574 144 591
rect 114 557 144 574
rect 114 540 121 557
rect 138 540 144 557
rect 114 523 144 540
rect 114 506 121 523
rect 138 506 144 523
rect 114 489 144 506
rect 114 472 121 489
rect 138 472 144 489
rect 114 455 144 472
rect 114 438 121 455
rect 138 438 144 455
rect 114 421 144 438
rect 114 404 121 421
rect 138 404 144 421
rect 114 387 144 404
rect 114 370 121 387
rect 138 370 144 387
rect 114 353 144 370
rect 114 336 121 353
rect 138 336 144 353
rect 114 319 144 336
rect 114 302 121 319
rect 138 302 144 319
rect 114 285 144 302
rect 114 268 121 285
rect 138 268 144 285
rect 114 251 144 268
rect 114 234 121 251
rect 138 234 144 251
rect 114 217 144 234
rect 114 200 121 217
rect 138 200 144 217
rect 114 183 144 200
rect 114 166 121 183
rect 138 166 144 183
rect 114 150 144 166
rect 159 1135 189 1150
rect 159 1118 165 1135
rect 182 1118 189 1135
rect 159 1101 189 1118
rect 159 1084 165 1101
rect 182 1084 189 1101
rect 159 1067 189 1084
rect 159 1050 165 1067
rect 182 1050 189 1067
rect 159 1033 189 1050
rect 159 1016 165 1033
rect 182 1016 189 1033
rect 159 999 189 1016
rect 159 982 166 999
rect 183 982 189 999
rect 159 965 189 982
rect 159 948 166 965
rect 183 948 189 965
rect 159 931 189 948
rect 159 914 166 931
rect 183 914 189 931
rect 159 897 189 914
rect 159 880 166 897
rect 183 880 189 897
rect 159 863 189 880
rect 159 846 166 863
rect 183 846 189 863
rect 159 829 189 846
rect 159 812 166 829
rect 183 812 189 829
rect 159 795 189 812
rect 159 778 166 795
rect 183 778 189 795
rect 159 761 189 778
rect 159 744 166 761
rect 183 744 189 761
rect 159 727 189 744
rect 159 710 166 727
rect 183 710 189 727
rect 159 693 189 710
rect 159 676 166 693
rect 183 676 189 693
rect 159 659 189 676
rect 159 642 166 659
rect 183 642 189 659
rect 159 625 189 642
rect 159 608 166 625
rect 183 608 189 625
rect 159 591 189 608
rect 159 574 166 591
rect 183 574 189 591
rect 159 557 189 574
rect 159 540 166 557
rect 183 540 189 557
rect 159 523 189 540
rect 159 506 166 523
rect 183 506 189 523
rect 159 489 189 506
rect 159 472 166 489
rect 183 472 189 489
rect 159 455 189 472
rect 159 438 166 455
rect 183 438 189 455
rect 159 421 189 438
rect 159 404 166 421
rect 183 404 189 421
rect 159 387 189 404
rect 159 370 166 387
rect 183 370 189 387
rect 159 353 189 370
rect 159 336 166 353
rect 183 336 189 353
rect 159 319 189 336
rect 159 302 166 319
rect 183 302 189 319
rect 159 285 189 302
rect 159 268 166 285
rect 183 268 189 285
rect 159 251 189 268
rect 159 234 166 251
rect 183 234 189 251
rect 159 217 189 234
rect 159 200 166 217
rect 183 200 189 217
rect 159 183 189 200
rect 159 166 166 183
rect 183 166 189 183
rect 159 150 189 166
rect 204 1135 234 1150
rect 204 1118 210 1135
rect 227 1118 234 1135
rect 204 1101 234 1118
rect 204 1084 210 1101
rect 227 1084 234 1101
rect 204 1067 234 1084
rect 204 1050 210 1067
rect 227 1050 234 1067
rect 204 1033 234 1050
rect 204 1016 210 1033
rect 227 1016 234 1033
rect 204 999 234 1016
rect 204 982 211 999
rect 228 982 234 999
rect 204 965 234 982
rect 204 948 211 965
rect 228 948 234 965
rect 204 931 234 948
rect 204 914 211 931
rect 228 914 234 931
rect 204 897 234 914
rect 204 880 211 897
rect 228 880 234 897
rect 204 863 234 880
rect 204 846 211 863
rect 228 846 234 863
rect 204 829 234 846
rect 204 812 211 829
rect 228 812 234 829
rect 204 795 234 812
rect 204 778 211 795
rect 228 778 234 795
rect 204 761 234 778
rect 204 744 211 761
rect 228 744 234 761
rect 204 727 234 744
rect 204 710 211 727
rect 228 710 234 727
rect 204 693 234 710
rect 204 676 211 693
rect 228 676 234 693
rect 204 659 234 676
rect 204 642 211 659
rect 228 642 234 659
rect 204 625 234 642
rect 204 608 211 625
rect 228 608 234 625
rect 204 591 234 608
rect 204 574 211 591
rect 228 574 234 591
rect 204 557 234 574
rect 204 540 211 557
rect 228 540 234 557
rect 204 523 234 540
rect 204 506 211 523
rect 228 506 234 523
rect 204 489 234 506
rect 204 472 211 489
rect 228 472 234 489
rect 204 455 234 472
rect 204 438 211 455
rect 228 438 234 455
rect 204 421 234 438
rect 204 404 211 421
rect 228 404 234 421
rect 204 387 234 404
rect 204 370 211 387
rect 228 370 234 387
rect 204 353 234 370
rect 204 336 211 353
rect 228 336 234 353
rect 204 319 234 336
rect 204 302 211 319
rect 228 302 234 319
rect 204 285 234 302
rect 204 268 211 285
rect 228 268 234 285
rect 204 251 234 268
rect 204 234 211 251
rect 228 234 234 251
rect 204 217 234 234
rect 204 200 211 217
rect 228 200 234 217
rect 204 183 234 200
rect 204 166 211 183
rect 228 166 234 183
rect 204 150 234 166
rect 249 1135 279 1150
rect 249 1118 255 1135
rect 272 1118 279 1135
rect 249 1101 279 1118
rect 249 1084 255 1101
rect 272 1084 279 1101
rect 249 1067 279 1084
rect 249 1050 255 1067
rect 272 1050 279 1067
rect 249 1033 279 1050
rect 249 1016 255 1033
rect 272 1016 279 1033
rect 249 999 279 1016
rect 249 982 256 999
rect 273 982 279 999
rect 249 965 279 982
rect 249 948 256 965
rect 273 948 279 965
rect 249 931 279 948
rect 249 914 256 931
rect 273 914 279 931
rect 249 897 279 914
rect 249 880 256 897
rect 273 880 279 897
rect 249 863 279 880
rect 249 846 256 863
rect 273 846 279 863
rect 249 829 279 846
rect 249 812 256 829
rect 273 812 279 829
rect 249 795 279 812
rect 249 778 256 795
rect 273 778 279 795
rect 249 761 279 778
rect 249 744 256 761
rect 273 744 279 761
rect 249 727 279 744
rect 249 710 256 727
rect 273 710 279 727
rect 249 693 279 710
rect 249 676 256 693
rect 273 676 279 693
rect 249 659 279 676
rect 249 642 256 659
rect 273 642 279 659
rect 249 625 279 642
rect 249 608 256 625
rect 273 608 279 625
rect 249 591 279 608
rect 249 574 256 591
rect 273 574 279 591
rect 249 557 279 574
rect 249 540 256 557
rect 273 540 279 557
rect 249 523 279 540
rect 249 506 256 523
rect 273 506 279 523
rect 249 489 279 506
rect 249 472 256 489
rect 273 472 279 489
rect 249 455 279 472
rect 249 438 256 455
rect 273 438 279 455
rect 249 421 279 438
rect 249 404 256 421
rect 273 404 279 421
rect 249 387 279 404
rect 249 370 256 387
rect 273 370 279 387
rect 249 353 279 370
rect 249 336 256 353
rect 273 336 279 353
rect 249 319 279 336
rect 249 302 256 319
rect 273 302 279 319
rect 249 285 279 302
rect 249 268 256 285
rect 273 268 279 285
rect 249 251 279 268
rect 249 234 256 251
rect 273 234 279 251
rect 249 217 279 234
rect 249 200 256 217
rect 273 200 279 217
rect 249 183 279 200
rect 249 166 256 183
rect 273 166 279 183
rect 249 150 279 166
rect 294 1135 325 1150
rect 294 1118 301 1135
rect 318 1118 325 1135
rect 294 1101 325 1118
rect 294 1084 301 1101
rect 318 1084 325 1101
rect 294 1067 325 1084
rect 294 1050 301 1067
rect 318 1050 325 1067
rect 294 1033 325 1050
rect 294 1016 301 1033
rect 318 1016 325 1033
rect 294 999 325 1016
rect 294 982 302 999
rect 319 982 325 999
rect 294 965 325 982
rect 294 948 302 965
rect 319 948 325 965
rect 294 931 325 948
rect 294 914 302 931
rect 319 914 325 931
rect 294 897 325 914
rect 294 880 302 897
rect 319 880 325 897
rect 294 863 325 880
rect 294 846 302 863
rect 319 846 325 863
rect 294 829 325 846
rect 294 812 302 829
rect 319 812 325 829
rect 294 795 325 812
rect 294 778 302 795
rect 319 778 325 795
rect 294 761 325 778
rect 294 744 302 761
rect 319 744 325 761
rect 294 727 325 744
rect 294 710 302 727
rect 319 710 325 727
rect 294 693 325 710
rect 294 676 302 693
rect 319 676 325 693
rect 294 659 325 676
rect 294 642 302 659
rect 319 642 325 659
rect 294 625 325 642
rect 294 608 302 625
rect 319 608 325 625
rect 294 591 325 608
rect 294 574 302 591
rect 319 574 325 591
rect 294 557 325 574
rect 294 540 302 557
rect 319 540 325 557
rect 294 523 325 540
rect 294 506 302 523
rect 319 506 325 523
rect 294 489 325 506
rect 294 472 302 489
rect 319 472 325 489
rect 294 455 325 472
rect 294 438 302 455
rect 319 438 325 455
rect 294 421 325 438
rect 294 404 302 421
rect 319 404 325 421
rect 294 387 325 404
rect 294 370 302 387
rect 319 370 325 387
rect 294 353 325 370
rect 294 336 302 353
rect 319 336 325 353
rect 294 319 325 336
rect 294 302 302 319
rect 319 302 325 319
rect 294 285 325 302
rect 294 268 302 285
rect 319 268 325 285
rect 294 251 325 268
rect 294 234 302 251
rect 319 234 325 251
rect 294 217 325 234
rect 294 200 302 217
rect 319 200 325 217
rect 294 183 325 200
rect 294 166 302 183
rect 319 166 325 183
rect 294 150 325 166
rect 340 1137 369 1150
rect 340 1120 346 1137
rect 363 1120 369 1137
rect 340 1103 369 1120
rect 340 1086 346 1103
rect 363 1086 369 1103
rect 340 1069 369 1086
rect 340 1052 346 1069
rect 363 1052 369 1069
rect 340 1035 369 1052
rect 340 1018 346 1035
rect 363 1018 369 1035
rect 340 1001 369 1018
rect 340 984 346 1001
rect 363 984 369 1001
rect 340 967 369 984
rect 340 950 346 967
rect 363 950 369 967
rect 340 933 369 950
rect 340 916 346 933
rect 363 916 369 933
rect 340 899 369 916
rect 340 882 346 899
rect 363 882 369 899
rect 340 865 369 882
rect 340 848 346 865
rect 363 848 369 865
rect 340 831 369 848
rect 340 814 346 831
rect 363 814 369 831
rect 340 797 369 814
rect 340 780 346 797
rect 363 780 369 797
rect 340 763 369 780
rect 340 746 346 763
rect 363 746 369 763
rect 340 729 369 746
rect 340 712 346 729
rect 363 712 369 729
rect 340 695 369 712
rect 340 678 346 695
rect 363 678 369 695
rect 340 661 369 678
rect 340 644 346 661
rect 363 644 369 661
rect 340 627 369 644
rect 340 610 346 627
rect 363 610 369 627
rect 340 593 369 610
rect 340 576 346 593
rect 363 576 369 593
rect 340 559 369 576
rect 340 542 346 559
rect 363 542 369 559
rect 340 525 369 542
rect 340 508 346 525
rect 363 508 369 525
rect 340 491 369 508
rect 340 474 346 491
rect 363 474 369 491
rect 340 457 369 474
rect 340 440 346 457
rect 363 440 369 457
rect 340 423 369 440
rect 340 406 346 423
rect 363 406 369 423
rect 340 389 369 406
rect 340 372 346 389
rect 363 372 369 389
rect 340 355 369 372
rect 340 338 346 355
rect 363 338 369 355
rect 340 321 369 338
rect 340 304 346 321
rect 363 304 369 321
rect 340 287 369 304
rect 340 270 346 287
rect 363 270 369 287
rect 340 253 369 270
rect 340 236 346 253
rect 363 236 369 253
rect 340 219 369 236
rect 340 202 346 219
rect 363 202 369 219
rect 340 185 369 202
rect 340 168 346 185
rect 363 168 369 185
rect 340 150 369 168
rect 384 1135 414 1150
rect 384 1118 390 1135
rect 407 1118 414 1135
rect 384 1101 414 1118
rect 384 1084 390 1101
rect 407 1084 414 1101
rect 384 1067 414 1084
rect 384 1050 390 1067
rect 407 1050 414 1067
rect 384 1033 414 1050
rect 384 1016 390 1033
rect 407 1016 414 1033
rect 384 999 414 1016
rect 384 982 391 999
rect 408 982 414 999
rect 384 965 414 982
rect 384 948 391 965
rect 408 948 414 965
rect 384 931 414 948
rect 384 914 391 931
rect 408 914 414 931
rect 384 897 414 914
rect 384 880 391 897
rect 408 880 414 897
rect 384 863 414 880
rect 384 846 391 863
rect 408 846 414 863
rect 384 829 414 846
rect 384 812 391 829
rect 408 812 414 829
rect 384 795 414 812
rect 384 778 391 795
rect 408 778 414 795
rect 384 761 414 778
rect 384 744 391 761
rect 408 744 414 761
rect 384 727 414 744
rect 384 710 391 727
rect 408 710 414 727
rect 384 693 414 710
rect 384 676 391 693
rect 408 676 414 693
rect 384 659 414 676
rect 384 642 391 659
rect 408 642 414 659
rect 384 625 414 642
rect 384 608 391 625
rect 408 608 414 625
rect 384 591 414 608
rect 384 574 391 591
rect 408 574 414 591
rect 384 557 414 574
rect 384 540 391 557
rect 408 540 414 557
rect 384 523 414 540
rect 384 506 391 523
rect 408 506 414 523
rect 384 489 414 506
rect 384 472 391 489
rect 408 472 414 489
rect 384 455 414 472
rect 384 438 391 455
rect 408 438 414 455
rect 384 421 414 438
rect 384 404 391 421
rect 408 404 414 421
rect 384 387 414 404
rect 384 370 391 387
rect 408 370 414 387
rect 384 353 414 370
rect 384 336 391 353
rect 408 336 414 353
rect 384 319 414 336
rect 384 302 391 319
rect 408 302 414 319
rect 384 285 414 302
rect 384 268 391 285
rect 408 268 414 285
rect 384 251 414 268
rect 384 234 391 251
rect 408 234 414 251
rect 384 217 414 234
rect 384 200 391 217
rect 408 200 414 217
rect 384 183 414 200
rect 384 166 391 183
rect 408 166 414 183
rect 384 150 414 166
rect 429 1135 459 1150
rect 429 1118 435 1135
rect 452 1118 459 1135
rect 429 1101 459 1118
rect 429 1084 435 1101
rect 452 1084 459 1101
rect 429 1067 459 1084
rect 429 1050 435 1067
rect 452 1050 459 1067
rect 429 1033 459 1050
rect 429 1016 435 1033
rect 452 1016 459 1033
rect 429 999 459 1016
rect 429 982 436 999
rect 453 982 459 999
rect 429 965 459 982
rect 429 948 436 965
rect 453 948 459 965
rect 429 931 459 948
rect 429 914 436 931
rect 453 914 459 931
rect 429 897 459 914
rect 429 880 436 897
rect 453 880 459 897
rect 429 863 459 880
rect 429 846 436 863
rect 453 846 459 863
rect 429 829 459 846
rect 429 812 436 829
rect 453 812 459 829
rect 429 795 459 812
rect 429 778 436 795
rect 453 778 459 795
rect 429 761 459 778
rect 429 744 436 761
rect 453 744 459 761
rect 429 727 459 744
rect 429 710 436 727
rect 453 710 459 727
rect 429 693 459 710
rect 429 676 436 693
rect 453 676 459 693
rect 429 659 459 676
rect 429 642 436 659
rect 453 642 459 659
rect 429 625 459 642
rect 429 608 436 625
rect 453 608 459 625
rect 429 591 459 608
rect 429 574 436 591
rect 453 574 459 591
rect 429 557 459 574
rect 429 540 436 557
rect 453 540 459 557
rect 429 523 459 540
rect 429 506 436 523
rect 453 506 459 523
rect 429 489 459 506
rect 429 472 436 489
rect 453 472 459 489
rect 429 455 459 472
rect 429 438 436 455
rect 453 438 459 455
rect 429 421 459 438
rect 429 404 436 421
rect 453 404 459 421
rect 429 387 459 404
rect 429 370 436 387
rect 453 370 459 387
rect 429 353 459 370
rect 429 336 436 353
rect 453 336 459 353
rect 429 319 459 336
rect 429 302 436 319
rect 453 302 459 319
rect 429 285 459 302
rect 429 268 436 285
rect 453 268 459 285
rect 429 251 459 268
rect 429 234 436 251
rect 453 234 459 251
rect 429 217 459 234
rect 429 200 436 217
rect 453 200 459 217
rect 429 183 459 200
rect 429 166 436 183
rect 453 166 459 183
rect 429 150 459 166
rect 474 1135 504 1150
rect 474 1118 480 1135
rect 497 1118 504 1135
rect 474 1101 504 1118
rect 474 1084 480 1101
rect 497 1084 504 1101
rect 474 1067 504 1084
rect 474 1050 480 1067
rect 497 1050 504 1067
rect 474 1033 504 1050
rect 474 1016 480 1033
rect 497 1016 504 1033
rect 474 999 504 1016
rect 474 982 481 999
rect 498 982 504 999
rect 474 965 504 982
rect 474 948 481 965
rect 498 948 504 965
rect 474 931 504 948
rect 474 914 481 931
rect 498 914 504 931
rect 474 897 504 914
rect 474 880 481 897
rect 498 880 504 897
rect 474 863 504 880
rect 474 846 481 863
rect 498 846 504 863
rect 474 829 504 846
rect 474 812 481 829
rect 498 812 504 829
rect 474 795 504 812
rect 474 778 481 795
rect 498 778 504 795
rect 474 761 504 778
rect 474 744 481 761
rect 498 744 504 761
rect 474 727 504 744
rect 474 710 481 727
rect 498 710 504 727
rect 474 693 504 710
rect 474 676 481 693
rect 498 676 504 693
rect 474 659 504 676
rect 474 642 481 659
rect 498 642 504 659
rect 474 625 504 642
rect 474 608 481 625
rect 498 608 504 625
rect 474 591 504 608
rect 474 574 481 591
rect 498 574 504 591
rect 474 557 504 574
rect 474 540 481 557
rect 498 540 504 557
rect 474 523 504 540
rect 474 506 481 523
rect 498 506 504 523
rect 474 489 504 506
rect 474 472 481 489
rect 498 472 504 489
rect 474 455 504 472
rect 474 438 481 455
rect 498 438 504 455
rect 474 421 504 438
rect 474 404 481 421
rect 498 404 504 421
rect 474 387 504 404
rect 474 370 481 387
rect 498 370 504 387
rect 474 353 504 370
rect 474 336 481 353
rect 498 336 504 353
rect 474 319 504 336
rect 474 302 481 319
rect 498 302 504 319
rect 474 285 504 302
rect 474 268 481 285
rect 498 268 504 285
rect 474 251 504 268
rect 474 234 481 251
rect 498 234 504 251
rect 474 217 504 234
rect 474 200 481 217
rect 498 200 504 217
rect 474 183 504 200
rect 474 166 481 183
rect 498 166 504 183
rect 474 150 504 166
rect 519 1135 549 1150
rect 519 1118 525 1135
rect 542 1118 549 1135
rect 519 1101 549 1118
rect 519 1084 525 1101
rect 542 1084 549 1101
rect 519 1067 549 1084
rect 519 1050 525 1067
rect 542 1050 549 1067
rect 519 1033 549 1050
rect 519 1016 525 1033
rect 542 1016 549 1033
rect 519 999 549 1016
rect 519 982 526 999
rect 543 982 549 999
rect 519 965 549 982
rect 519 948 526 965
rect 543 948 549 965
rect 519 931 549 948
rect 519 914 526 931
rect 543 914 549 931
rect 519 897 549 914
rect 519 880 526 897
rect 543 880 549 897
rect 519 863 549 880
rect 519 846 526 863
rect 543 846 549 863
rect 519 829 549 846
rect 519 812 526 829
rect 543 812 549 829
rect 519 795 549 812
rect 519 778 526 795
rect 543 778 549 795
rect 519 761 549 778
rect 519 744 526 761
rect 543 744 549 761
rect 519 727 549 744
rect 519 710 526 727
rect 543 710 549 727
rect 519 693 549 710
rect 519 676 526 693
rect 543 676 549 693
rect 519 659 549 676
rect 519 642 526 659
rect 543 642 549 659
rect 519 625 549 642
rect 519 608 526 625
rect 543 608 549 625
rect 519 591 549 608
rect 519 574 526 591
rect 543 574 549 591
rect 519 557 549 574
rect 519 540 526 557
rect 543 540 549 557
rect 519 523 549 540
rect 519 506 526 523
rect 543 506 549 523
rect 519 489 549 506
rect 519 472 526 489
rect 543 472 549 489
rect 519 455 549 472
rect 519 438 526 455
rect 543 438 549 455
rect 519 421 549 438
rect 519 404 526 421
rect 543 404 549 421
rect 519 387 549 404
rect 519 370 526 387
rect 543 370 549 387
rect 519 353 549 370
rect 519 336 526 353
rect 543 336 549 353
rect 519 319 549 336
rect 519 302 526 319
rect 543 302 549 319
rect 519 285 549 302
rect 519 268 526 285
rect 543 268 549 285
rect 519 251 549 268
rect 519 234 526 251
rect 543 234 549 251
rect 519 217 549 234
rect 519 200 526 217
rect 543 200 549 217
rect 519 183 549 200
rect 519 166 526 183
rect 543 166 549 183
rect 519 150 549 166
rect 564 1135 594 1150
rect 564 1118 570 1135
rect 587 1118 594 1135
rect 564 1101 594 1118
rect 564 1084 570 1101
rect 587 1084 594 1101
rect 564 1067 594 1084
rect 564 1050 570 1067
rect 587 1050 594 1067
rect 564 1033 594 1050
rect 564 1016 570 1033
rect 587 1016 594 1033
rect 564 999 594 1016
rect 564 982 571 999
rect 588 982 594 999
rect 564 965 594 982
rect 564 948 571 965
rect 588 948 594 965
rect 564 931 594 948
rect 564 914 571 931
rect 588 914 594 931
rect 564 897 594 914
rect 564 880 571 897
rect 588 880 594 897
rect 564 863 594 880
rect 564 846 571 863
rect 588 846 594 863
rect 564 829 594 846
rect 564 812 571 829
rect 588 812 594 829
rect 564 795 594 812
rect 564 778 571 795
rect 588 778 594 795
rect 564 761 594 778
rect 564 744 571 761
rect 588 744 594 761
rect 564 727 594 744
rect 564 710 571 727
rect 588 710 594 727
rect 564 693 594 710
rect 564 676 571 693
rect 588 676 594 693
rect 564 659 594 676
rect 564 642 571 659
rect 588 642 594 659
rect 564 625 594 642
rect 564 608 571 625
rect 588 608 594 625
rect 564 591 594 608
rect 564 574 571 591
rect 588 574 594 591
rect 564 557 594 574
rect 564 540 571 557
rect 588 540 594 557
rect 564 523 594 540
rect 564 506 571 523
rect 588 506 594 523
rect 564 489 594 506
rect 564 472 571 489
rect 588 472 594 489
rect 564 455 594 472
rect 564 438 571 455
rect 588 438 594 455
rect 564 421 594 438
rect 564 404 571 421
rect 588 404 594 421
rect 564 387 594 404
rect 564 370 571 387
rect 588 370 594 387
rect 564 353 594 370
rect 564 336 571 353
rect 588 336 594 353
rect 564 319 594 336
rect 564 302 571 319
rect 588 302 594 319
rect 564 285 594 302
rect 564 268 571 285
rect 588 268 594 285
rect 564 251 594 268
rect 564 234 571 251
rect 588 234 594 251
rect 564 217 594 234
rect 564 200 571 217
rect 588 200 594 217
rect 564 183 594 200
rect 564 166 571 183
rect 588 166 594 183
rect 564 150 594 166
rect 609 1135 639 1150
rect 609 1118 615 1135
rect 632 1118 639 1135
rect 609 1101 639 1118
rect 609 1084 615 1101
rect 632 1084 639 1101
rect 609 1067 639 1084
rect 609 1050 615 1067
rect 632 1050 639 1067
rect 609 1033 639 1050
rect 609 1016 615 1033
rect 632 1016 639 1033
rect 609 999 639 1016
rect 609 982 616 999
rect 633 982 639 999
rect 609 965 639 982
rect 609 948 616 965
rect 633 948 639 965
rect 609 931 639 948
rect 609 914 616 931
rect 633 914 639 931
rect 609 897 639 914
rect 609 880 616 897
rect 633 880 639 897
rect 609 863 639 880
rect 609 846 616 863
rect 633 846 639 863
rect 609 829 639 846
rect 609 812 616 829
rect 633 812 639 829
rect 609 795 639 812
rect 609 778 616 795
rect 633 778 639 795
rect 609 761 639 778
rect 609 744 616 761
rect 633 744 639 761
rect 609 727 639 744
rect 609 710 616 727
rect 633 710 639 727
rect 609 693 639 710
rect 609 676 616 693
rect 633 676 639 693
rect 609 659 639 676
rect 609 642 616 659
rect 633 642 639 659
rect 609 625 639 642
rect 609 608 616 625
rect 633 608 639 625
rect 609 591 639 608
rect 609 574 616 591
rect 633 574 639 591
rect 609 557 639 574
rect 609 540 616 557
rect 633 540 639 557
rect 609 523 639 540
rect 609 506 616 523
rect 633 506 639 523
rect 609 489 639 506
rect 609 472 616 489
rect 633 472 639 489
rect 609 455 639 472
rect 609 438 616 455
rect 633 438 639 455
rect 609 421 639 438
rect 609 404 616 421
rect 633 404 639 421
rect 609 387 639 404
rect 609 370 616 387
rect 633 370 639 387
rect 609 353 639 370
rect 609 336 616 353
rect 633 336 639 353
rect 609 319 639 336
rect 609 302 616 319
rect 633 302 639 319
rect 609 285 639 302
rect 609 268 616 285
rect 633 268 639 285
rect 609 251 639 268
rect 609 234 616 251
rect 633 234 639 251
rect 609 217 639 234
rect 609 200 616 217
rect 633 200 639 217
rect 609 183 639 200
rect 609 166 616 183
rect 633 166 639 183
rect 609 150 639 166
rect 654 1135 684 1150
rect 654 1118 660 1135
rect 677 1118 684 1135
rect 654 1101 684 1118
rect 654 1084 660 1101
rect 677 1084 684 1101
rect 654 1067 684 1084
rect 654 1050 660 1067
rect 677 1050 684 1067
rect 654 1033 684 1050
rect 654 1016 660 1033
rect 677 1016 684 1033
rect 654 999 684 1016
rect 654 982 661 999
rect 678 982 684 999
rect 654 965 684 982
rect 654 948 661 965
rect 678 948 684 965
rect 654 931 684 948
rect 654 914 661 931
rect 678 914 684 931
rect 654 897 684 914
rect 654 880 661 897
rect 678 880 684 897
rect 654 863 684 880
rect 654 846 661 863
rect 678 846 684 863
rect 654 829 684 846
rect 654 812 661 829
rect 678 812 684 829
rect 654 795 684 812
rect 654 778 661 795
rect 678 778 684 795
rect 654 761 684 778
rect 654 744 661 761
rect 678 744 684 761
rect 654 727 684 744
rect 654 710 661 727
rect 678 710 684 727
rect 654 693 684 710
rect 654 676 661 693
rect 678 676 684 693
rect 654 659 684 676
rect 654 642 661 659
rect 678 642 684 659
rect 654 625 684 642
rect 654 608 661 625
rect 678 608 684 625
rect 654 591 684 608
rect 654 574 661 591
rect 678 574 684 591
rect 654 557 684 574
rect 654 540 661 557
rect 678 540 684 557
rect 654 523 684 540
rect 654 506 661 523
rect 678 506 684 523
rect 654 489 684 506
rect 654 472 661 489
rect 678 472 684 489
rect 654 455 684 472
rect 654 438 661 455
rect 678 438 684 455
rect 654 421 684 438
rect 654 404 661 421
rect 678 404 684 421
rect 654 387 684 404
rect 654 370 661 387
rect 678 370 684 387
rect 654 353 684 370
rect 654 336 661 353
rect 678 336 684 353
rect 654 319 684 336
rect 654 302 661 319
rect 678 302 684 319
rect 654 285 684 302
rect 654 268 661 285
rect 678 268 684 285
rect 654 251 684 268
rect 654 234 661 251
rect 678 234 684 251
rect 654 217 684 234
rect 654 200 661 217
rect 678 200 684 217
rect 654 183 684 200
rect 654 166 661 183
rect 678 166 684 183
rect 654 150 684 166
rect 699 1137 728 1150
rect 699 1120 705 1137
rect 722 1120 728 1137
rect 699 1103 728 1120
rect 699 1086 705 1103
rect 722 1086 728 1103
rect 699 1069 728 1086
rect 699 1052 705 1069
rect 722 1052 728 1069
rect 699 1035 728 1052
rect 699 1018 705 1035
rect 722 1018 728 1035
rect 699 1001 728 1018
rect 699 984 705 1001
rect 722 984 728 1001
rect 699 967 728 984
rect 699 950 705 967
rect 722 950 728 967
rect 699 933 728 950
rect 699 916 705 933
rect 722 916 728 933
rect 699 899 728 916
rect 699 882 705 899
rect 722 882 728 899
rect 699 865 728 882
rect 699 848 705 865
rect 722 848 728 865
rect 699 831 728 848
rect 699 814 705 831
rect 722 814 728 831
rect 699 797 728 814
rect 699 780 705 797
rect 722 780 728 797
rect 699 763 728 780
rect 699 746 705 763
rect 722 746 728 763
rect 699 729 728 746
rect 699 712 705 729
rect 722 712 728 729
rect 699 695 728 712
rect 699 678 705 695
rect 722 678 728 695
rect 699 661 728 678
rect 699 644 705 661
rect 722 644 728 661
rect 699 627 728 644
rect 699 610 705 627
rect 722 610 728 627
rect 699 593 728 610
rect 699 576 705 593
rect 722 576 728 593
rect 699 559 728 576
rect 699 542 705 559
rect 722 542 728 559
rect 699 525 728 542
rect 699 508 705 525
rect 722 508 728 525
rect 699 491 728 508
rect 699 474 705 491
rect 722 474 728 491
rect 699 457 728 474
rect 699 440 705 457
rect 722 440 728 457
rect 699 423 728 440
rect 699 406 705 423
rect 722 406 728 423
rect 699 389 728 406
rect 699 372 705 389
rect 722 372 728 389
rect 699 355 728 372
rect 699 338 705 355
rect 722 338 728 355
rect 699 321 728 338
rect 699 304 705 321
rect 722 304 728 321
rect 699 287 728 304
rect 699 270 705 287
rect 722 270 728 287
rect 699 253 728 270
rect 699 236 705 253
rect 722 236 728 253
rect 699 219 728 236
rect 699 202 705 219
rect 722 202 728 219
rect 699 185 728 202
rect 699 168 705 185
rect 722 168 728 185
rect 699 150 728 168
rect 743 1135 773 1150
rect 743 1118 749 1135
rect 766 1118 773 1135
rect 743 1101 773 1118
rect 743 1084 749 1101
rect 766 1084 773 1101
rect 743 1067 773 1084
rect 743 1050 749 1067
rect 766 1050 773 1067
rect 743 1033 773 1050
rect 743 1016 749 1033
rect 766 1016 773 1033
rect 743 999 773 1016
rect 743 982 750 999
rect 767 982 773 999
rect 743 965 773 982
rect 743 948 750 965
rect 767 948 773 965
rect 743 931 773 948
rect 743 914 750 931
rect 767 914 773 931
rect 743 897 773 914
rect 743 880 750 897
rect 767 880 773 897
rect 743 863 773 880
rect 743 846 750 863
rect 767 846 773 863
rect 743 829 773 846
rect 743 812 750 829
rect 767 812 773 829
rect 743 795 773 812
rect 743 778 750 795
rect 767 778 773 795
rect 743 761 773 778
rect 743 744 750 761
rect 767 744 773 761
rect 743 727 773 744
rect 743 710 750 727
rect 767 710 773 727
rect 743 693 773 710
rect 743 676 750 693
rect 767 676 773 693
rect 743 659 773 676
rect 743 642 750 659
rect 767 642 773 659
rect 743 625 773 642
rect 743 608 750 625
rect 767 608 773 625
rect 743 591 773 608
rect 743 574 750 591
rect 767 574 773 591
rect 743 557 773 574
rect 743 540 750 557
rect 767 540 773 557
rect 743 523 773 540
rect 743 506 750 523
rect 767 506 773 523
rect 743 489 773 506
rect 743 472 750 489
rect 767 472 773 489
rect 743 455 773 472
rect 743 438 750 455
rect 767 438 773 455
rect 743 421 773 438
rect 743 404 750 421
rect 767 404 773 421
rect 743 387 773 404
rect 743 370 750 387
rect 767 370 773 387
rect 743 353 773 370
rect 743 336 750 353
rect 767 336 773 353
rect 743 319 773 336
rect 743 302 750 319
rect 767 302 773 319
rect 743 285 773 302
rect 743 268 750 285
rect 767 268 773 285
rect 743 251 773 268
rect 743 234 750 251
rect 767 234 773 251
rect 743 217 773 234
rect 743 200 750 217
rect 767 200 773 217
rect 743 183 773 200
rect 743 166 750 183
rect 767 166 773 183
rect 743 150 773 166
rect 788 1135 818 1150
rect 788 1118 794 1135
rect 811 1118 818 1135
rect 788 1101 818 1118
rect 788 1084 794 1101
rect 811 1084 818 1101
rect 788 1067 818 1084
rect 788 1050 794 1067
rect 811 1050 818 1067
rect 788 1033 818 1050
rect 788 1016 794 1033
rect 811 1016 818 1033
rect 788 999 818 1016
rect 788 982 795 999
rect 812 982 818 999
rect 788 965 818 982
rect 788 948 795 965
rect 812 948 818 965
rect 788 931 818 948
rect 788 914 795 931
rect 812 914 818 931
rect 788 897 818 914
rect 788 880 795 897
rect 812 880 818 897
rect 788 863 818 880
rect 788 846 795 863
rect 812 846 818 863
rect 788 829 818 846
rect 788 812 795 829
rect 812 812 818 829
rect 788 795 818 812
rect 788 778 795 795
rect 812 778 818 795
rect 788 761 818 778
rect 788 744 795 761
rect 812 744 818 761
rect 788 727 818 744
rect 788 710 795 727
rect 812 710 818 727
rect 788 693 818 710
rect 788 676 795 693
rect 812 676 818 693
rect 788 659 818 676
rect 788 642 795 659
rect 812 642 818 659
rect 788 625 818 642
rect 788 608 795 625
rect 812 608 818 625
rect 788 591 818 608
rect 788 574 795 591
rect 812 574 818 591
rect 788 557 818 574
rect 788 540 795 557
rect 812 540 818 557
rect 788 523 818 540
rect 788 506 795 523
rect 812 506 818 523
rect 788 489 818 506
rect 788 472 795 489
rect 812 472 818 489
rect 788 455 818 472
rect 788 438 795 455
rect 812 438 818 455
rect 788 421 818 438
rect 788 404 795 421
rect 812 404 818 421
rect 788 387 818 404
rect 788 370 795 387
rect 812 370 818 387
rect 788 353 818 370
rect 788 336 795 353
rect 812 336 818 353
rect 788 319 818 336
rect 788 302 795 319
rect 812 302 818 319
rect 788 285 818 302
rect 788 268 795 285
rect 812 268 818 285
rect 788 251 818 268
rect 788 234 795 251
rect 812 234 818 251
rect 788 217 818 234
rect 788 200 795 217
rect 812 200 818 217
rect 788 183 818 200
rect 788 166 795 183
rect 812 166 818 183
rect 788 150 818 166
rect 833 1135 863 1150
rect 833 1118 839 1135
rect 856 1118 863 1135
rect 833 1101 863 1118
rect 833 1084 839 1101
rect 856 1084 863 1101
rect 833 1067 863 1084
rect 833 1050 839 1067
rect 856 1050 863 1067
rect 833 1033 863 1050
rect 833 1016 839 1033
rect 856 1016 863 1033
rect 833 999 863 1016
rect 833 982 840 999
rect 857 982 863 999
rect 833 965 863 982
rect 833 948 840 965
rect 857 948 863 965
rect 833 931 863 948
rect 833 914 840 931
rect 857 914 863 931
rect 833 897 863 914
rect 833 880 840 897
rect 857 880 863 897
rect 833 863 863 880
rect 833 846 840 863
rect 857 846 863 863
rect 833 829 863 846
rect 833 812 840 829
rect 857 812 863 829
rect 833 795 863 812
rect 833 778 840 795
rect 857 778 863 795
rect 833 761 863 778
rect 833 744 840 761
rect 857 744 863 761
rect 833 727 863 744
rect 833 710 840 727
rect 857 710 863 727
rect 833 693 863 710
rect 833 676 840 693
rect 857 676 863 693
rect 833 659 863 676
rect 833 642 840 659
rect 857 642 863 659
rect 833 625 863 642
rect 833 608 840 625
rect 857 608 863 625
rect 833 591 863 608
rect 833 574 840 591
rect 857 574 863 591
rect 833 557 863 574
rect 833 540 840 557
rect 857 540 863 557
rect 833 523 863 540
rect 833 506 840 523
rect 857 506 863 523
rect 833 489 863 506
rect 833 472 840 489
rect 857 472 863 489
rect 833 455 863 472
rect 833 438 840 455
rect 857 438 863 455
rect 833 421 863 438
rect 833 404 840 421
rect 857 404 863 421
rect 833 387 863 404
rect 833 370 840 387
rect 857 370 863 387
rect 833 353 863 370
rect 833 336 840 353
rect 857 336 863 353
rect 833 319 863 336
rect 833 302 840 319
rect 857 302 863 319
rect 833 285 863 302
rect 833 268 840 285
rect 857 268 863 285
rect 833 251 863 268
rect 833 234 840 251
rect 857 234 863 251
rect 833 217 863 234
rect 833 200 840 217
rect 857 200 863 217
rect 833 183 863 200
rect 833 166 840 183
rect 857 166 863 183
rect 833 150 863 166
rect 878 1135 908 1150
rect 878 1118 884 1135
rect 901 1118 908 1135
rect 878 1101 908 1118
rect 878 1084 884 1101
rect 901 1084 908 1101
rect 878 1067 908 1084
rect 878 1050 884 1067
rect 901 1050 908 1067
rect 878 1033 908 1050
rect 878 1016 884 1033
rect 901 1016 908 1033
rect 878 999 908 1016
rect 878 982 885 999
rect 902 982 908 999
rect 878 965 908 982
rect 878 948 885 965
rect 902 948 908 965
rect 878 931 908 948
rect 878 914 885 931
rect 902 914 908 931
rect 878 897 908 914
rect 878 880 885 897
rect 902 880 908 897
rect 878 863 908 880
rect 878 846 885 863
rect 902 846 908 863
rect 878 829 908 846
rect 878 812 885 829
rect 902 812 908 829
rect 878 795 908 812
rect 878 778 885 795
rect 902 778 908 795
rect 878 761 908 778
rect 878 744 885 761
rect 902 744 908 761
rect 878 727 908 744
rect 878 710 885 727
rect 902 710 908 727
rect 878 693 908 710
rect 878 676 885 693
rect 902 676 908 693
rect 878 659 908 676
rect 878 642 885 659
rect 902 642 908 659
rect 878 625 908 642
rect 878 608 885 625
rect 902 608 908 625
rect 878 591 908 608
rect 878 574 885 591
rect 902 574 908 591
rect 878 557 908 574
rect 878 540 885 557
rect 902 540 908 557
rect 878 523 908 540
rect 878 506 885 523
rect 902 506 908 523
rect 878 489 908 506
rect 878 472 885 489
rect 902 472 908 489
rect 878 455 908 472
rect 878 438 885 455
rect 902 438 908 455
rect 878 421 908 438
rect 878 404 885 421
rect 902 404 908 421
rect 878 387 908 404
rect 878 370 885 387
rect 902 370 908 387
rect 878 353 908 370
rect 878 336 885 353
rect 902 336 908 353
rect 878 319 908 336
rect 878 302 885 319
rect 902 302 908 319
rect 878 285 908 302
rect 878 268 885 285
rect 902 268 908 285
rect 878 251 908 268
rect 878 234 885 251
rect 902 234 908 251
rect 878 217 908 234
rect 878 200 885 217
rect 902 200 908 217
rect 878 183 908 200
rect 878 166 885 183
rect 902 166 908 183
rect 878 150 908 166
rect 923 1135 953 1150
rect 923 1118 929 1135
rect 946 1118 953 1135
rect 923 1101 953 1118
rect 923 1084 929 1101
rect 946 1084 953 1101
rect 923 1067 953 1084
rect 923 1050 929 1067
rect 946 1050 953 1067
rect 923 1033 953 1050
rect 923 1016 929 1033
rect 946 1016 953 1033
rect 923 999 953 1016
rect 923 982 930 999
rect 947 982 953 999
rect 923 965 953 982
rect 923 948 930 965
rect 947 948 953 965
rect 923 931 953 948
rect 923 914 930 931
rect 947 914 953 931
rect 923 897 953 914
rect 923 880 930 897
rect 947 880 953 897
rect 923 863 953 880
rect 923 846 930 863
rect 947 846 953 863
rect 923 829 953 846
rect 923 812 930 829
rect 947 812 953 829
rect 923 795 953 812
rect 923 778 930 795
rect 947 778 953 795
rect 923 761 953 778
rect 923 744 930 761
rect 947 744 953 761
rect 923 727 953 744
rect 923 710 930 727
rect 947 710 953 727
rect 923 693 953 710
rect 923 676 930 693
rect 947 676 953 693
rect 923 659 953 676
rect 923 642 930 659
rect 947 642 953 659
rect 923 625 953 642
rect 923 608 930 625
rect 947 608 953 625
rect 923 591 953 608
rect 923 574 930 591
rect 947 574 953 591
rect 923 557 953 574
rect 923 540 930 557
rect 947 540 953 557
rect 923 523 953 540
rect 923 506 930 523
rect 947 506 953 523
rect 923 489 953 506
rect 923 472 930 489
rect 947 472 953 489
rect 923 455 953 472
rect 923 438 930 455
rect 947 438 953 455
rect 923 421 953 438
rect 923 404 930 421
rect 947 404 953 421
rect 923 387 953 404
rect 923 370 930 387
rect 947 370 953 387
rect 923 353 953 370
rect 923 336 930 353
rect 947 336 953 353
rect 923 319 953 336
rect 923 302 930 319
rect 947 302 953 319
rect 923 285 953 302
rect 923 268 930 285
rect 947 268 953 285
rect 923 251 953 268
rect 923 234 930 251
rect 947 234 953 251
rect 923 217 953 234
rect 923 200 930 217
rect 947 200 953 217
rect 923 183 953 200
rect 923 166 930 183
rect 947 166 953 183
rect 923 150 953 166
rect 968 1135 998 1150
rect 968 1118 974 1135
rect 991 1118 998 1135
rect 968 1101 998 1118
rect 968 1084 974 1101
rect 991 1084 998 1101
rect 968 1067 998 1084
rect 968 1050 974 1067
rect 991 1050 998 1067
rect 968 1033 998 1050
rect 968 1016 974 1033
rect 991 1016 998 1033
rect 968 999 998 1016
rect 968 982 975 999
rect 992 982 998 999
rect 968 965 998 982
rect 968 948 975 965
rect 992 948 998 965
rect 968 931 998 948
rect 968 914 975 931
rect 992 914 998 931
rect 968 897 998 914
rect 968 880 975 897
rect 992 880 998 897
rect 968 863 998 880
rect 968 846 975 863
rect 992 846 998 863
rect 968 829 998 846
rect 968 812 975 829
rect 992 812 998 829
rect 968 795 998 812
rect 968 778 975 795
rect 992 778 998 795
rect 968 761 998 778
rect 968 744 975 761
rect 992 744 998 761
rect 968 727 998 744
rect 968 710 975 727
rect 992 710 998 727
rect 968 693 998 710
rect 968 676 975 693
rect 992 676 998 693
rect 968 659 998 676
rect 968 642 975 659
rect 992 642 998 659
rect 968 625 998 642
rect 968 608 975 625
rect 992 608 998 625
rect 968 591 998 608
rect 968 574 975 591
rect 992 574 998 591
rect 968 557 998 574
rect 968 540 975 557
rect 992 540 998 557
rect 968 523 998 540
rect 968 506 975 523
rect 992 506 998 523
rect 968 489 998 506
rect 968 472 975 489
rect 992 472 998 489
rect 968 455 998 472
rect 968 438 975 455
rect 992 438 998 455
rect 968 421 998 438
rect 968 404 975 421
rect 992 404 998 421
rect 968 387 998 404
rect 968 370 975 387
rect 992 370 998 387
rect 968 353 998 370
rect 968 336 975 353
rect 992 336 998 353
rect 968 319 998 336
rect 968 302 975 319
rect 992 302 998 319
rect 968 285 998 302
rect 968 268 975 285
rect 992 268 998 285
rect 968 251 998 268
rect 968 234 975 251
rect 992 234 998 251
rect 968 217 998 234
rect 968 200 975 217
rect 992 200 998 217
rect 968 183 998 200
rect 968 166 975 183
rect 992 166 998 183
rect 968 150 998 166
rect 1013 1135 1044 1150
rect 1013 1118 1020 1135
rect 1037 1118 1044 1135
rect 1013 1101 1044 1118
rect 1013 1084 1020 1101
rect 1037 1084 1044 1101
rect 1013 1067 1044 1084
rect 1013 1050 1020 1067
rect 1037 1050 1044 1067
rect 1013 1033 1044 1050
rect 1013 1016 1020 1033
rect 1037 1016 1044 1033
rect 1013 999 1044 1016
rect 1013 982 1021 999
rect 1038 982 1044 999
rect 1013 965 1044 982
rect 1013 948 1021 965
rect 1038 948 1044 965
rect 1013 931 1044 948
rect 1013 914 1021 931
rect 1038 914 1044 931
rect 1013 897 1044 914
rect 1013 880 1021 897
rect 1038 880 1044 897
rect 1013 863 1044 880
rect 1013 846 1021 863
rect 1038 846 1044 863
rect 1013 829 1044 846
rect 1013 812 1021 829
rect 1038 812 1044 829
rect 1013 795 1044 812
rect 1013 778 1021 795
rect 1038 778 1044 795
rect 1013 761 1044 778
rect 1013 744 1021 761
rect 1038 744 1044 761
rect 1013 727 1044 744
rect 1013 710 1021 727
rect 1038 710 1044 727
rect 1013 693 1044 710
rect 1013 676 1021 693
rect 1038 676 1044 693
rect 1013 659 1044 676
rect 1013 642 1021 659
rect 1038 642 1044 659
rect 1013 625 1044 642
rect 1013 608 1021 625
rect 1038 608 1044 625
rect 1013 591 1044 608
rect 1013 574 1021 591
rect 1038 574 1044 591
rect 1013 557 1044 574
rect 1013 540 1021 557
rect 1038 540 1044 557
rect 1013 523 1044 540
rect 1013 506 1021 523
rect 1038 506 1044 523
rect 1013 489 1044 506
rect 1013 472 1021 489
rect 1038 472 1044 489
rect 1013 455 1044 472
rect 1013 438 1021 455
rect 1038 438 1044 455
rect 1013 421 1044 438
rect 1013 404 1021 421
rect 1038 404 1044 421
rect 1013 387 1044 404
rect 1013 370 1021 387
rect 1038 370 1044 387
rect 1013 353 1044 370
rect 1013 336 1021 353
rect 1038 336 1044 353
rect 1013 319 1044 336
rect 1013 302 1021 319
rect 1038 302 1044 319
rect 1013 285 1044 302
rect 1013 268 1021 285
rect 1038 268 1044 285
rect 1013 251 1044 268
rect 1013 234 1021 251
rect 1038 234 1044 251
rect 1013 217 1044 234
rect 1013 200 1021 217
rect 1038 200 1044 217
rect 1013 183 1044 200
rect 1013 166 1021 183
rect 1038 166 1044 183
rect 1013 150 1044 166
rect 1059 1137 1088 1150
rect 1059 1120 1065 1137
rect 1082 1120 1088 1137
rect 1059 1103 1088 1120
rect 1059 1086 1065 1103
rect 1082 1086 1088 1103
rect 1059 1069 1088 1086
rect 1059 1052 1065 1069
rect 1082 1052 1088 1069
rect 1059 1035 1088 1052
rect 1059 1018 1065 1035
rect 1082 1018 1088 1035
rect 1059 1001 1088 1018
rect 1059 984 1065 1001
rect 1082 984 1088 1001
rect 1059 967 1088 984
rect 1059 950 1065 967
rect 1082 950 1088 967
rect 1059 933 1088 950
rect 1059 916 1065 933
rect 1082 916 1088 933
rect 1059 899 1088 916
rect 1059 882 1065 899
rect 1082 882 1088 899
rect 1059 865 1088 882
rect 1059 848 1065 865
rect 1082 848 1088 865
rect 1059 831 1088 848
rect 1059 814 1065 831
rect 1082 814 1088 831
rect 1059 797 1088 814
rect 1059 780 1065 797
rect 1082 780 1088 797
rect 1059 763 1088 780
rect 1059 746 1065 763
rect 1082 746 1088 763
rect 1059 729 1088 746
rect 1059 712 1065 729
rect 1082 712 1088 729
rect 1059 695 1088 712
rect 1059 678 1065 695
rect 1082 678 1088 695
rect 1059 661 1088 678
rect 1059 644 1065 661
rect 1082 644 1088 661
rect 1059 627 1088 644
rect 1059 610 1065 627
rect 1082 610 1088 627
rect 1059 593 1088 610
rect 1059 576 1065 593
rect 1082 576 1088 593
rect 1059 559 1088 576
rect 1059 542 1065 559
rect 1082 542 1088 559
rect 1059 525 1088 542
rect 1059 508 1065 525
rect 1082 508 1088 525
rect 1059 491 1088 508
rect 1059 474 1065 491
rect 1082 474 1088 491
rect 1059 457 1088 474
rect 1059 440 1065 457
rect 1082 440 1088 457
rect 1059 423 1088 440
rect 1059 406 1065 423
rect 1082 406 1088 423
rect 1059 389 1088 406
rect 1059 372 1065 389
rect 1082 372 1088 389
rect 1059 355 1088 372
rect 1059 338 1065 355
rect 1082 338 1088 355
rect 1059 321 1088 338
rect 1059 304 1065 321
rect 1082 304 1088 321
rect 1059 287 1088 304
rect 1059 270 1065 287
rect 1082 270 1088 287
rect 1059 253 1088 270
rect 1059 236 1065 253
rect 1082 236 1088 253
rect 1059 219 1088 236
rect 1059 202 1065 219
rect 1082 202 1088 219
rect 1059 185 1088 202
rect 1059 168 1065 185
rect 1082 168 1088 185
rect 1059 150 1088 168
rect 1103 1135 1133 1150
rect 1103 1118 1109 1135
rect 1126 1118 1133 1135
rect 1103 1101 1133 1118
rect 1103 1084 1109 1101
rect 1126 1084 1133 1101
rect 1103 1067 1133 1084
rect 1103 1050 1109 1067
rect 1126 1050 1133 1067
rect 1103 1033 1133 1050
rect 1103 1016 1109 1033
rect 1126 1016 1133 1033
rect 1103 999 1133 1016
rect 1103 982 1110 999
rect 1127 982 1133 999
rect 1103 965 1133 982
rect 1103 948 1110 965
rect 1127 948 1133 965
rect 1103 931 1133 948
rect 1103 914 1110 931
rect 1127 914 1133 931
rect 1103 897 1133 914
rect 1103 880 1110 897
rect 1127 880 1133 897
rect 1103 863 1133 880
rect 1103 846 1110 863
rect 1127 846 1133 863
rect 1103 829 1133 846
rect 1103 812 1110 829
rect 1127 812 1133 829
rect 1103 795 1133 812
rect 1103 778 1110 795
rect 1127 778 1133 795
rect 1103 761 1133 778
rect 1103 744 1110 761
rect 1127 744 1133 761
rect 1103 727 1133 744
rect 1103 710 1110 727
rect 1127 710 1133 727
rect 1103 693 1133 710
rect 1103 676 1110 693
rect 1127 676 1133 693
rect 1103 659 1133 676
rect 1103 642 1110 659
rect 1127 642 1133 659
rect 1103 625 1133 642
rect 1103 608 1110 625
rect 1127 608 1133 625
rect 1103 591 1133 608
rect 1103 574 1110 591
rect 1127 574 1133 591
rect 1103 557 1133 574
rect 1103 540 1110 557
rect 1127 540 1133 557
rect 1103 523 1133 540
rect 1103 506 1110 523
rect 1127 506 1133 523
rect 1103 489 1133 506
rect 1103 472 1110 489
rect 1127 472 1133 489
rect 1103 455 1133 472
rect 1103 438 1110 455
rect 1127 438 1133 455
rect 1103 421 1133 438
rect 1103 404 1110 421
rect 1127 404 1133 421
rect 1103 387 1133 404
rect 1103 370 1110 387
rect 1127 370 1133 387
rect 1103 353 1133 370
rect 1103 336 1110 353
rect 1127 336 1133 353
rect 1103 319 1133 336
rect 1103 302 1110 319
rect 1127 302 1133 319
rect 1103 285 1133 302
rect 1103 268 1110 285
rect 1127 268 1133 285
rect 1103 251 1133 268
rect 1103 234 1110 251
rect 1127 234 1133 251
rect 1103 217 1133 234
rect 1103 200 1110 217
rect 1127 200 1133 217
rect 1103 183 1133 200
rect 1103 166 1110 183
rect 1127 166 1133 183
rect 1103 150 1133 166
rect 1148 1135 1178 1150
rect 1148 1118 1154 1135
rect 1171 1118 1178 1135
rect 1148 1101 1178 1118
rect 1148 1084 1154 1101
rect 1171 1084 1178 1101
rect 1148 1067 1178 1084
rect 1148 1050 1154 1067
rect 1171 1050 1178 1067
rect 1148 1033 1178 1050
rect 1148 1016 1154 1033
rect 1171 1016 1178 1033
rect 1148 999 1178 1016
rect 1148 982 1155 999
rect 1172 982 1178 999
rect 1148 965 1178 982
rect 1148 948 1155 965
rect 1172 948 1178 965
rect 1148 931 1178 948
rect 1148 914 1155 931
rect 1172 914 1178 931
rect 1148 897 1178 914
rect 1148 880 1155 897
rect 1172 880 1178 897
rect 1148 863 1178 880
rect 1148 846 1155 863
rect 1172 846 1178 863
rect 1148 829 1178 846
rect 1148 812 1155 829
rect 1172 812 1178 829
rect 1148 795 1178 812
rect 1148 778 1155 795
rect 1172 778 1178 795
rect 1148 761 1178 778
rect 1148 744 1155 761
rect 1172 744 1178 761
rect 1148 727 1178 744
rect 1148 710 1155 727
rect 1172 710 1178 727
rect 1148 693 1178 710
rect 1148 676 1155 693
rect 1172 676 1178 693
rect 1148 659 1178 676
rect 1148 642 1155 659
rect 1172 642 1178 659
rect 1148 625 1178 642
rect 1148 608 1155 625
rect 1172 608 1178 625
rect 1148 591 1178 608
rect 1148 574 1155 591
rect 1172 574 1178 591
rect 1148 557 1178 574
rect 1148 540 1155 557
rect 1172 540 1178 557
rect 1148 523 1178 540
rect 1148 506 1155 523
rect 1172 506 1178 523
rect 1148 489 1178 506
rect 1148 472 1155 489
rect 1172 472 1178 489
rect 1148 455 1178 472
rect 1148 438 1155 455
rect 1172 438 1178 455
rect 1148 421 1178 438
rect 1148 404 1155 421
rect 1172 404 1178 421
rect 1148 387 1178 404
rect 1148 370 1155 387
rect 1172 370 1178 387
rect 1148 353 1178 370
rect 1148 336 1155 353
rect 1172 336 1178 353
rect 1148 319 1178 336
rect 1148 302 1155 319
rect 1172 302 1178 319
rect 1148 285 1178 302
rect 1148 268 1155 285
rect 1172 268 1178 285
rect 1148 251 1178 268
rect 1148 234 1155 251
rect 1172 234 1178 251
rect 1148 217 1178 234
rect 1148 200 1155 217
rect 1172 200 1178 217
rect 1148 183 1178 200
rect 1148 166 1155 183
rect 1172 166 1178 183
rect 1148 150 1178 166
rect 1193 1135 1223 1150
rect 1193 1118 1199 1135
rect 1216 1118 1223 1135
rect 1193 1101 1223 1118
rect 1193 1084 1199 1101
rect 1216 1084 1223 1101
rect 1193 1067 1223 1084
rect 1193 1050 1199 1067
rect 1216 1050 1223 1067
rect 1193 1033 1223 1050
rect 1193 1016 1199 1033
rect 1216 1016 1223 1033
rect 1193 999 1223 1016
rect 1193 982 1200 999
rect 1217 982 1223 999
rect 1193 965 1223 982
rect 1193 948 1200 965
rect 1217 948 1223 965
rect 1193 931 1223 948
rect 1193 914 1200 931
rect 1217 914 1223 931
rect 1193 897 1223 914
rect 1193 880 1200 897
rect 1217 880 1223 897
rect 1193 863 1223 880
rect 1193 846 1200 863
rect 1217 846 1223 863
rect 1193 829 1223 846
rect 1193 812 1200 829
rect 1217 812 1223 829
rect 1193 795 1223 812
rect 1193 778 1200 795
rect 1217 778 1223 795
rect 1193 761 1223 778
rect 1193 744 1200 761
rect 1217 744 1223 761
rect 1193 727 1223 744
rect 1193 710 1200 727
rect 1217 710 1223 727
rect 1193 693 1223 710
rect 1193 676 1200 693
rect 1217 676 1223 693
rect 1193 659 1223 676
rect 1193 642 1200 659
rect 1217 642 1223 659
rect 1193 625 1223 642
rect 1193 608 1200 625
rect 1217 608 1223 625
rect 1193 591 1223 608
rect 1193 574 1200 591
rect 1217 574 1223 591
rect 1193 557 1223 574
rect 1193 540 1200 557
rect 1217 540 1223 557
rect 1193 523 1223 540
rect 1193 506 1200 523
rect 1217 506 1223 523
rect 1193 489 1223 506
rect 1193 472 1200 489
rect 1217 472 1223 489
rect 1193 455 1223 472
rect 1193 438 1200 455
rect 1217 438 1223 455
rect 1193 421 1223 438
rect 1193 404 1200 421
rect 1217 404 1223 421
rect 1193 387 1223 404
rect 1193 370 1200 387
rect 1217 370 1223 387
rect 1193 353 1223 370
rect 1193 336 1200 353
rect 1217 336 1223 353
rect 1193 319 1223 336
rect 1193 302 1200 319
rect 1217 302 1223 319
rect 1193 285 1223 302
rect 1193 268 1200 285
rect 1217 268 1223 285
rect 1193 251 1223 268
rect 1193 234 1200 251
rect 1217 234 1223 251
rect 1193 217 1223 234
rect 1193 200 1200 217
rect 1217 200 1223 217
rect 1193 183 1223 200
rect 1193 166 1200 183
rect 1217 166 1223 183
rect 1193 150 1223 166
rect 1238 1135 1268 1150
rect 1238 1118 1244 1135
rect 1261 1118 1268 1135
rect 1238 1101 1268 1118
rect 1238 1084 1244 1101
rect 1261 1084 1268 1101
rect 1238 1067 1268 1084
rect 1238 1050 1244 1067
rect 1261 1050 1268 1067
rect 1238 1033 1268 1050
rect 1238 1016 1244 1033
rect 1261 1016 1268 1033
rect 1238 999 1268 1016
rect 1238 982 1245 999
rect 1262 982 1268 999
rect 1238 965 1268 982
rect 1238 948 1245 965
rect 1262 948 1268 965
rect 1238 931 1268 948
rect 1238 914 1245 931
rect 1262 914 1268 931
rect 1238 897 1268 914
rect 1238 880 1245 897
rect 1262 880 1268 897
rect 1238 863 1268 880
rect 1238 846 1245 863
rect 1262 846 1268 863
rect 1238 829 1268 846
rect 1238 812 1245 829
rect 1262 812 1268 829
rect 1238 795 1268 812
rect 1238 778 1245 795
rect 1262 778 1268 795
rect 1238 761 1268 778
rect 1238 744 1245 761
rect 1262 744 1268 761
rect 1238 727 1268 744
rect 1238 710 1245 727
rect 1262 710 1268 727
rect 1238 693 1268 710
rect 1238 676 1245 693
rect 1262 676 1268 693
rect 1238 659 1268 676
rect 1238 642 1245 659
rect 1262 642 1268 659
rect 1238 625 1268 642
rect 1238 608 1245 625
rect 1262 608 1268 625
rect 1238 591 1268 608
rect 1238 574 1245 591
rect 1262 574 1268 591
rect 1238 557 1268 574
rect 1238 540 1245 557
rect 1262 540 1268 557
rect 1238 523 1268 540
rect 1238 506 1245 523
rect 1262 506 1268 523
rect 1238 489 1268 506
rect 1238 472 1245 489
rect 1262 472 1268 489
rect 1238 455 1268 472
rect 1238 438 1245 455
rect 1262 438 1268 455
rect 1238 421 1268 438
rect 1238 404 1245 421
rect 1262 404 1268 421
rect 1238 387 1268 404
rect 1238 370 1245 387
rect 1262 370 1268 387
rect 1238 353 1268 370
rect 1238 336 1245 353
rect 1262 336 1268 353
rect 1238 319 1268 336
rect 1238 302 1245 319
rect 1262 302 1268 319
rect 1238 285 1268 302
rect 1238 268 1245 285
rect 1262 268 1268 285
rect 1238 251 1268 268
rect 1238 234 1245 251
rect 1262 234 1268 251
rect 1238 217 1268 234
rect 1238 200 1245 217
rect 1262 200 1268 217
rect 1238 183 1268 200
rect 1238 166 1245 183
rect 1262 166 1268 183
rect 1238 150 1268 166
rect 1283 1135 1313 1150
rect 1283 1118 1289 1135
rect 1306 1118 1313 1135
rect 1283 1101 1313 1118
rect 1283 1084 1289 1101
rect 1306 1084 1313 1101
rect 1283 1067 1313 1084
rect 1283 1050 1289 1067
rect 1306 1050 1313 1067
rect 1283 1033 1313 1050
rect 1283 1016 1289 1033
rect 1306 1016 1313 1033
rect 1283 999 1313 1016
rect 1283 982 1290 999
rect 1307 982 1313 999
rect 1283 965 1313 982
rect 1283 948 1290 965
rect 1307 948 1313 965
rect 1283 931 1313 948
rect 1283 914 1290 931
rect 1307 914 1313 931
rect 1283 897 1313 914
rect 1283 880 1290 897
rect 1307 880 1313 897
rect 1283 863 1313 880
rect 1283 846 1290 863
rect 1307 846 1313 863
rect 1283 829 1313 846
rect 1283 812 1290 829
rect 1307 812 1313 829
rect 1283 795 1313 812
rect 1283 778 1290 795
rect 1307 778 1313 795
rect 1283 761 1313 778
rect 1283 744 1290 761
rect 1307 744 1313 761
rect 1283 727 1313 744
rect 1283 710 1290 727
rect 1307 710 1313 727
rect 1283 693 1313 710
rect 1283 676 1290 693
rect 1307 676 1313 693
rect 1283 659 1313 676
rect 1283 642 1290 659
rect 1307 642 1313 659
rect 1283 625 1313 642
rect 1283 608 1290 625
rect 1307 608 1313 625
rect 1283 591 1313 608
rect 1283 574 1290 591
rect 1307 574 1313 591
rect 1283 557 1313 574
rect 1283 540 1290 557
rect 1307 540 1313 557
rect 1283 523 1313 540
rect 1283 506 1290 523
rect 1307 506 1313 523
rect 1283 489 1313 506
rect 1283 472 1290 489
rect 1307 472 1313 489
rect 1283 455 1313 472
rect 1283 438 1290 455
rect 1307 438 1313 455
rect 1283 421 1313 438
rect 1283 404 1290 421
rect 1307 404 1313 421
rect 1283 387 1313 404
rect 1283 370 1290 387
rect 1307 370 1313 387
rect 1283 353 1313 370
rect 1283 336 1290 353
rect 1307 336 1313 353
rect 1283 319 1313 336
rect 1283 302 1290 319
rect 1307 302 1313 319
rect 1283 285 1313 302
rect 1283 268 1290 285
rect 1307 268 1313 285
rect 1283 251 1313 268
rect 1283 234 1290 251
rect 1307 234 1313 251
rect 1283 217 1313 234
rect 1283 200 1290 217
rect 1307 200 1313 217
rect 1283 183 1313 200
rect 1283 166 1290 183
rect 1307 166 1313 183
rect 1283 150 1313 166
rect 1328 1135 1358 1150
rect 1328 1118 1334 1135
rect 1351 1118 1358 1135
rect 1328 1101 1358 1118
rect 1328 1084 1334 1101
rect 1351 1084 1358 1101
rect 1328 1067 1358 1084
rect 1328 1050 1334 1067
rect 1351 1050 1358 1067
rect 1328 1033 1358 1050
rect 1328 1016 1334 1033
rect 1351 1016 1358 1033
rect 1328 999 1358 1016
rect 1328 982 1335 999
rect 1352 982 1358 999
rect 1328 965 1358 982
rect 1328 948 1335 965
rect 1352 948 1358 965
rect 1328 931 1358 948
rect 1328 914 1335 931
rect 1352 914 1358 931
rect 1328 897 1358 914
rect 1328 880 1335 897
rect 1352 880 1358 897
rect 1328 863 1358 880
rect 1328 846 1335 863
rect 1352 846 1358 863
rect 1328 829 1358 846
rect 1328 812 1335 829
rect 1352 812 1358 829
rect 1328 795 1358 812
rect 1328 778 1335 795
rect 1352 778 1358 795
rect 1328 761 1358 778
rect 1328 744 1335 761
rect 1352 744 1358 761
rect 1328 727 1358 744
rect 1328 710 1335 727
rect 1352 710 1358 727
rect 1328 693 1358 710
rect 1328 676 1335 693
rect 1352 676 1358 693
rect 1328 659 1358 676
rect 1328 642 1335 659
rect 1352 642 1358 659
rect 1328 625 1358 642
rect 1328 608 1335 625
rect 1352 608 1358 625
rect 1328 591 1358 608
rect 1328 574 1335 591
rect 1352 574 1358 591
rect 1328 557 1358 574
rect 1328 540 1335 557
rect 1352 540 1358 557
rect 1328 523 1358 540
rect 1328 506 1335 523
rect 1352 506 1358 523
rect 1328 489 1358 506
rect 1328 472 1335 489
rect 1352 472 1358 489
rect 1328 455 1358 472
rect 1328 438 1335 455
rect 1352 438 1358 455
rect 1328 421 1358 438
rect 1328 404 1335 421
rect 1352 404 1358 421
rect 1328 387 1358 404
rect 1328 370 1335 387
rect 1352 370 1358 387
rect 1328 353 1358 370
rect 1328 336 1335 353
rect 1352 336 1358 353
rect 1328 319 1358 336
rect 1328 302 1335 319
rect 1352 302 1358 319
rect 1328 285 1358 302
rect 1328 268 1335 285
rect 1352 268 1358 285
rect 1328 251 1358 268
rect 1328 234 1335 251
rect 1352 234 1358 251
rect 1328 217 1358 234
rect 1328 200 1335 217
rect 1352 200 1358 217
rect 1328 183 1358 200
rect 1328 166 1335 183
rect 1352 166 1358 183
rect 1328 150 1358 166
rect 1373 1135 1403 1150
rect 1373 1118 1379 1135
rect 1396 1118 1403 1135
rect 1373 1101 1403 1118
rect 1373 1084 1379 1101
rect 1396 1084 1403 1101
rect 1373 1067 1403 1084
rect 1373 1050 1379 1067
rect 1396 1050 1403 1067
rect 1373 1033 1403 1050
rect 1373 1016 1379 1033
rect 1396 1016 1403 1033
rect 1373 999 1403 1016
rect 1373 982 1380 999
rect 1397 982 1403 999
rect 1373 965 1403 982
rect 1373 948 1380 965
rect 1397 948 1403 965
rect 1373 931 1403 948
rect 1373 914 1380 931
rect 1397 914 1403 931
rect 1373 897 1403 914
rect 1373 880 1380 897
rect 1397 880 1403 897
rect 1373 863 1403 880
rect 1373 846 1380 863
rect 1397 846 1403 863
rect 1373 829 1403 846
rect 1373 812 1380 829
rect 1397 812 1403 829
rect 1373 795 1403 812
rect 1373 778 1380 795
rect 1397 778 1403 795
rect 1373 761 1403 778
rect 1373 744 1380 761
rect 1397 744 1403 761
rect 1373 727 1403 744
rect 1373 710 1380 727
rect 1397 710 1403 727
rect 1373 693 1403 710
rect 1373 676 1380 693
rect 1397 676 1403 693
rect 1373 659 1403 676
rect 1373 642 1380 659
rect 1397 642 1403 659
rect 1373 625 1403 642
rect 1373 608 1380 625
rect 1397 608 1403 625
rect 1373 591 1403 608
rect 1373 574 1380 591
rect 1397 574 1403 591
rect 1373 557 1403 574
rect 1373 540 1380 557
rect 1397 540 1403 557
rect 1373 523 1403 540
rect 1373 506 1380 523
rect 1397 506 1403 523
rect 1373 489 1403 506
rect 1373 472 1380 489
rect 1397 472 1403 489
rect 1373 455 1403 472
rect 1373 438 1380 455
rect 1397 438 1403 455
rect 1373 421 1403 438
rect 1373 404 1380 421
rect 1397 404 1403 421
rect 1373 387 1403 404
rect 1373 370 1380 387
rect 1397 370 1403 387
rect 1373 353 1403 370
rect 1373 336 1380 353
rect 1397 336 1403 353
rect 1373 319 1403 336
rect 1373 302 1380 319
rect 1397 302 1403 319
rect 1373 285 1403 302
rect 1373 268 1380 285
rect 1397 268 1403 285
rect 1373 251 1403 268
rect 1373 234 1380 251
rect 1397 234 1403 251
rect 1373 217 1403 234
rect 1373 200 1380 217
rect 1397 200 1403 217
rect 1373 183 1403 200
rect 1373 166 1380 183
rect 1397 166 1403 183
rect 1373 150 1403 166
rect 1418 1137 1447 1150
rect 1418 1120 1424 1137
rect 1441 1120 1447 1137
rect 1418 1103 1447 1120
rect 1418 1086 1424 1103
rect 1441 1086 1447 1103
rect 1418 1069 1447 1086
rect 1418 1052 1424 1069
rect 1441 1052 1447 1069
rect 1418 1035 1447 1052
rect 1418 1018 1424 1035
rect 1441 1018 1447 1035
rect 1418 1001 1447 1018
rect 1418 984 1424 1001
rect 1441 984 1447 1001
rect 1418 967 1447 984
rect 1418 950 1424 967
rect 1441 950 1447 967
rect 1418 933 1447 950
rect 1418 916 1424 933
rect 1441 916 1447 933
rect 1418 899 1447 916
rect 1418 882 1424 899
rect 1441 882 1447 899
rect 1418 865 1447 882
rect 1418 848 1424 865
rect 1441 848 1447 865
rect 1418 831 1447 848
rect 1418 814 1424 831
rect 1441 814 1447 831
rect 1418 797 1447 814
rect 1418 780 1424 797
rect 1441 780 1447 797
rect 1418 763 1447 780
rect 1418 746 1424 763
rect 1441 746 1447 763
rect 1418 729 1447 746
rect 1418 712 1424 729
rect 1441 712 1447 729
rect 1418 695 1447 712
rect 1418 678 1424 695
rect 1441 678 1447 695
rect 1418 661 1447 678
rect 1418 644 1424 661
rect 1441 644 1447 661
rect 1418 627 1447 644
rect 1418 610 1424 627
rect 1441 610 1447 627
rect 1418 593 1447 610
rect 1418 576 1424 593
rect 1441 576 1447 593
rect 1418 559 1447 576
rect 1418 542 1424 559
rect 1441 542 1447 559
rect 1418 525 1447 542
rect 1418 508 1424 525
rect 1441 508 1447 525
rect 1418 491 1447 508
rect 1418 474 1424 491
rect 1441 474 1447 491
rect 1418 457 1447 474
rect 1418 440 1424 457
rect 1441 440 1447 457
rect 1418 423 1447 440
rect 1418 406 1424 423
rect 1441 406 1447 423
rect 1418 389 1447 406
rect 1418 372 1424 389
rect 1441 372 1447 389
rect 1418 355 1447 372
rect 1418 338 1424 355
rect 1441 338 1447 355
rect 1418 321 1447 338
rect 1418 304 1424 321
rect 1441 304 1447 321
rect 1418 287 1447 304
rect 1418 270 1424 287
rect 1441 270 1447 287
rect 1418 253 1447 270
rect 1418 236 1424 253
rect 1441 236 1447 253
rect 1418 219 1447 236
rect 1418 202 1424 219
rect 1441 202 1447 219
rect 1418 185 1447 202
rect 1418 168 1424 185
rect 1441 168 1447 185
rect 1418 150 1447 168
rect 1462 1135 1492 1150
rect 1462 1118 1468 1135
rect 1485 1118 1492 1135
rect 1462 1101 1492 1118
rect 1462 1084 1468 1101
rect 1485 1084 1492 1101
rect 1462 1067 1492 1084
rect 1462 1050 1468 1067
rect 1485 1050 1492 1067
rect 1462 1033 1492 1050
rect 1462 1016 1468 1033
rect 1485 1016 1492 1033
rect 1462 999 1492 1016
rect 1462 982 1469 999
rect 1486 982 1492 999
rect 1462 965 1492 982
rect 1462 948 1469 965
rect 1486 948 1492 965
rect 1462 931 1492 948
rect 1462 914 1469 931
rect 1486 914 1492 931
rect 1462 897 1492 914
rect 1462 880 1469 897
rect 1486 880 1492 897
rect 1462 863 1492 880
rect 1462 846 1469 863
rect 1486 846 1492 863
rect 1462 829 1492 846
rect 1462 812 1469 829
rect 1486 812 1492 829
rect 1462 795 1492 812
rect 1462 778 1469 795
rect 1486 778 1492 795
rect 1462 761 1492 778
rect 1462 744 1469 761
rect 1486 744 1492 761
rect 1462 727 1492 744
rect 1462 710 1469 727
rect 1486 710 1492 727
rect 1462 693 1492 710
rect 1462 676 1469 693
rect 1486 676 1492 693
rect 1462 659 1492 676
rect 1462 642 1469 659
rect 1486 642 1492 659
rect 1462 625 1492 642
rect 1462 608 1469 625
rect 1486 608 1492 625
rect 1462 591 1492 608
rect 1462 574 1469 591
rect 1486 574 1492 591
rect 1462 557 1492 574
rect 1462 540 1469 557
rect 1486 540 1492 557
rect 1462 523 1492 540
rect 1462 506 1469 523
rect 1486 506 1492 523
rect 1462 489 1492 506
rect 1462 472 1469 489
rect 1486 472 1492 489
rect 1462 455 1492 472
rect 1462 438 1469 455
rect 1486 438 1492 455
rect 1462 421 1492 438
rect 1462 404 1469 421
rect 1486 404 1492 421
rect 1462 387 1492 404
rect 1462 370 1469 387
rect 1486 370 1492 387
rect 1462 353 1492 370
rect 1462 336 1469 353
rect 1486 336 1492 353
rect 1462 319 1492 336
rect 1462 302 1469 319
rect 1486 302 1492 319
rect 1462 285 1492 302
rect 1462 268 1469 285
rect 1486 268 1492 285
rect 1462 251 1492 268
rect 1462 234 1469 251
rect 1486 234 1492 251
rect 1462 217 1492 234
rect 1462 200 1469 217
rect 1486 200 1492 217
rect 1462 183 1492 200
rect 1462 166 1469 183
rect 1486 166 1492 183
rect 1462 150 1492 166
rect 1507 1135 1537 1150
rect 1507 1118 1513 1135
rect 1530 1118 1537 1135
rect 1507 1101 1537 1118
rect 1507 1084 1513 1101
rect 1530 1084 1537 1101
rect 1507 1067 1537 1084
rect 1507 1050 1513 1067
rect 1530 1050 1537 1067
rect 1507 1033 1537 1050
rect 1507 1016 1513 1033
rect 1530 1016 1537 1033
rect 1507 999 1537 1016
rect 1507 982 1514 999
rect 1531 982 1537 999
rect 1507 965 1537 982
rect 1507 948 1514 965
rect 1531 948 1537 965
rect 1507 931 1537 948
rect 1507 914 1514 931
rect 1531 914 1537 931
rect 1507 897 1537 914
rect 1507 880 1514 897
rect 1531 880 1537 897
rect 1507 863 1537 880
rect 1507 846 1514 863
rect 1531 846 1537 863
rect 1507 829 1537 846
rect 1507 812 1514 829
rect 1531 812 1537 829
rect 1507 795 1537 812
rect 1507 778 1514 795
rect 1531 778 1537 795
rect 1507 761 1537 778
rect 1507 744 1514 761
rect 1531 744 1537 761
rect 1507 727 1537 744
rect 1507 710 1514 727
rect 1531 710 1537 727
rect 1507 693 1537 710
rect 1507 676 1514 693
rect 1531 676 1537 693
rect 1507 659 1537 676
rect 1507 642 1514 659
rect 1531 642 1537 659
rect 1507 625 1537 642
rect 1507 608 1514 625
rect 1531 608 1537 625
rect 1507 591 1537 608
rect 1507 574 1514 591
rect 1531 574 1537 591
rect 1507 557 1537 574
rect 1507 540 1514 557
rect 1531 540 1537 557
rect 1507 523 1537 540
rect 1507 506 1514 523
rect 1531 506 1537 523
rect 1507 489 1537 506
rect 1507 472 1514 489
rect 1531 472 1537 489
rect 1507 455 1537 472
rect 1507 438 1514 455
rect 1531 438 1537 455
rect 1507 421 1537 438
rect 1507 404 1514 421
rect 1531 404 1537 421
rect 1507 387 1537 404
rect 1507 370 1514 387
rect 1531 370 1537 387
rect 1507 353 1537 370
rect 1507 336 1514 353
rect 1531 336 1537 353
rect 1507 319 1537 336
rect 1507 302 1514 319
rect 1531 302 1537 319
rect 1507 285 1537 302
rect 1507 268 1514 285
rect 1531 268 1537 285
rect 1507 251 1537 268
rect 1507 234 1514 251
rect 1531 234 1537 251
rect 1507 217 1537 234
rect 1507 200 1514 217
rect 1531 200 1537 217
rect 1507 183 1537 200
rect 1507 166 1514 183
rect 1531 166 1537 183
rect 1507 150 1537 166
rect 1552 1135 1582 1150
rect 1552 1118 1558 1135
rect 1575 1118 1582 1135
rect 1552 1101 1582 1118
rect 1552 1084 1558 1101
rect 1575 1084 1582 1101
rect 1552 1067 1582 1084
rect 1552 1050 1558 1067
rect 1575 1050 1582 1067
rect 1552 1033 1582 1050
rect 1552 1016 1558 1033
rect 1575 1016 1582 1033
rect 1552 999 1582 1016
rect 1552 982 1559 999
rect 1576 982 1582 999
rect 1552 965 1582 982
rect 1552 948 1559 965
rect 1576 948 1582 965
rect 1552 931 1582 948
rect 1552 914 1559 931
rect 1576 914 1582 931
rect 1552 897 1582 914
rect 1552 880 1559 897
rect 1576 880 1582 897
rect 1552 863 1582 880
rect 1552 846 1559 863
rect 1576 846 1582 863
rect 1552 829 1582 846
rect 1552 812 1559 829
rect 1576 812 1582 829
rect 1552 795 1582 812
rect 1552 778 1559 795
rect 1576 778 1582 795
rect 1552 761 1582 778
rect 1552 744 1559 761
rect 1576 744 1582 761
rect 1552 727 1582 744
rect 1552 710 1559 727
rect 1576 710 1582 727
rect 1552 693 1582 710
rect 1552 676 1559 693
rect 1576 676 1582 693
rect 1552 659 1582 676
rect 1552 642 1559 659
rect 1576 642 1582 659
rect 1552 625 1582 642
rect 1552 608 1559 625
rect 1576 608 1582 625
rect 1552 591 1582 608
rect 1552 574 1559 591
rect 1576 574 1582 591
rect 1552 557 1582 574
rect 1552 540 1559 557
rect 1576 540 1582 557
rect 1552 523 1582 540
rect 1552 506 1559 523
rect 1576 506 1582 523
rect 1552 489 1582 506
rect 1552 472 1559 489
rect 1576 472 1582 489
rect 1552 455 1582 472
rect 1552 438 1559 455
rect 1576 438 1582 455
rect 1552 421 1582 438
rect 1552 404 1559 421
rect 1576 404 1582 421
rect 1552 387 1582 404
rect 1552 370 1559 387
rect 1576 370 1582 387
rect 1552 353 1582 370
rect 1552 336 1559 353
rect 1576 336 1582 353
rect 1552 319 1582 336
rect 1552 302 1559 319
rect 1576 302 1582 319
rect 1552 285 1582 302
rect 1552 268 1559 285
rect 1576 268 1582 285
rect 1552 251 1582 268
rect 1552 234 1559 251
rect 1576 234 1582 251
rect 1552 217 1582 234
rect 1552 200 1559 217
rect 1576 200 1582 217
rect 1552 183 1582 200
rect 1552 166 1559 183
rect 1576 166 1582 183
rect 1552 150 1582 166
rect 1597 1135 1627 1150
rect 1597 1118 1603 1135
rect 1620 1118 1627 1135
rect 1597 1101 1627 1118
rect 1597 1084 1603 1101
rect 1620 1084 1627 1101
rect 1597 1067 1627 1084
rect 1597 1050 1603 1067
rect 1620 1050 1627 1067
rect 1597 1033 1627 1050
rect 1597 1016 1603 1033
rect 1620 1016 1627 1033
rect 1597 999 1627 1016
rect 1597 982 1604 999
rect 1621 982 1627 999
rect 1597 965 1627 982
rect 1597 948 1604 965
rect 1621 948 1627 965
rect 1597 931 1627 948
rect 1597 914 1604 931
rect 1621 914 1627 931
rect 1597 897 1627 914
rect 1597 880 1604 897
rect 1621 880 1627 897
rect 1597 863 1627 880
rect 1597 846 1604 863
rect 1621 846 1627 863
rect 1597 829 1627 846
rect 1597 812 1604 829
rect 1621 812 1627 829
rect 1597 795 1627 812
rect 1597 778 1604 795
rect 1621 778 1627 795
rect 1597 761 1627 778
rect 1597 744 1604 761
rect 1621 744 1627 761
rect 1597 727 1627 744
rect 1597 710 1604 727
rect 1621 710 1627 727
rect 1597 693 1627 710
rect 1597 676 1604 693
rect 1621 676 1627 693
rect 1597 659 1627 676
rect 1597 642 1604 659
rect 1621 642 1627 659
rect 1597 625 1627 642
rect 1597 608 1604 625
rect 1621 608 1627 625
rect 1597 591 1627 608
rect 1597 574 1604 591
rect 1621 574 1627 591
rect 1597 557 1627 574
rect 1597 540 1604 557
rect 1621 540 1627 557
rect 1597 523 1627 540
rect 1597 506 1604 523
rect 1621 506 1627 523
rect 1597 489 1627 506
rect 1597 472 1604 489
rect 1621 472 1627 489
rect 1597 455 1627 472
rect 1597 438 1604 455
rect 1621 438 1627 455
rect 1597 421 1627 438
rect 1597 404 1604 421
rect 1621 404 1627 421
rect 1597 387 1627 404
rect 1597 370 1604 387
rect 1621 370 1627 387
rect 1597 353 1627 370
rect 1597 336 1604 353
rect 1621 336 1627 353
rect 1597 319 1627 336
rect 1597 302 1604 319
rect 1621 302 1627 319
rect 1597 285 1627 302
rect 1597 268 1604 285
rect 1621 268 1627 285
rect 1597 251 1627 268
rect 1597 234 1604 251
rect 1621 234 1627 251
rect 1597 217 1627 234
rect 1597 200 1604 217
rect 1621 200 1627 217
rect 1597 183 1627 200
rect 1597 166 1604 183
rect 1621 166 1627 183
rect 1597 150 1627 166
rect 1642 1135 1672 1150
rect 1642 1118 1648 1135
rect 1665 1118 1672 1135
rect 1642 1101 1672 1118
rect 1642 1084 1648 1101
rect 1665 1084 1672 1101
rect 1642 1067 1672 1084
rect 1642 1050 1648 1067
rect 1665 1050 1672 1067
rect 1642 1033 1672 1050
rect 1642 1016 1648 1033
rect 1665 1016 1672 1033
rect 1642 999 1672 1016
rect 1642 982 1649 999
rect 1666 982 1672 999
rect 1642 965 1672 982
rect 1642 948 1649 965
rect 1666 948 1672 965
rect 1642 931 1672 948
rect 1642 914 1649 931
rect 1666 914 1672 931
rect 1642 897 1672 914
rect 1642 880 1649 897
rect 1666 880 1672 897
rect 1642 863 1672 880
rect 1642 846 1649 863
rect 1666 846 1672 863
rect 1642 829 1672 846
rect 1642 812 1649 829
rect 1666 812 1672 829
rect 1642 795 1672 812
rect 1642 778 1649 795
rect 1666 778 1672 795
rect 1642 761 1672 778
rect 1642 744 1649 761
rect 1666 744 1672 761
rect 1642 727 1672 744
rect 1642 710 1649 727
rect 1666 710 1672 727
rect 1642 693 1672 710
rect 1642 676 1649 693
rect 1666 676 1672 693
rect 1642 659 1672 676
rect 1642 642 1649 659
rect 1666 642 1672 659
rect 1642 625 1672 642
rect 1642 608 1649 625
rect 1666 608 1672 625
rect 1642 591 1672 608
rect 1642 574 1649 591
rect 1666 574 1672 591
rect 1642 557 1672 574
rect 1642 540 1649 557
rect 1666 540 1672 557
rect 1642 523 1672 540
rect 1642 506 1649 523
rect 1666 506 1672 523
rect 1642 489 1672 506
rect 1642 472 1649 489
rect 1666 472 1672 489
rect 1642 455 1672 472
rect 1642 438 1649 455
rect 1666 438 1672 455
rect 1642 421 1672 438
rect 1642 404 1649 421
rect 1666 404 1672 421
rect 1642 387 1672 404
rect 1642 370 1649 387
rect 1666 370 1672 387
rect 1642 353 1672 370
rect 1642 336 1649 353
rect 1666 336 1672 353
rect 1642 319 1672 336
rect 1642 302 1649 319
rect 1666 302 1672 319
rect 1642 285 1672 302
rect 1642 268 1649 285
rect 1666 268 1672 285
rect 1642 251 1672 268
rect 1642 234 1649 251
rect 1666 234 1672 251
rect 1642 217 1672 234
rect 1642 200 1649 217
rect 1666 200 1672 217
rect 1642 183 1672 200
rect 1642 166 1649 183
rect 1666 166 1672 183
rect 1642 150 1672 166
rect 1687 1135 1717 1150
rect 1687 1118 1693 1135
rect 1710 1118 1717 1135
rect 1687 1101 1717 1118
rect 1687 1084 1693 1101
rect 1710 1084 1717 1101
rect 1687 1067 1717 1084
rect 1687 1050 1693 1067
rect 1710 1050 1717 1067
rect 1687 1033 1717 1050
rect 1687 1016 1693 1033
rect 1710 1016 1717 1033
rect 1687 999 1717 1016
rect 1687 982 1694 999
rect 1711 982 1717 999
rect 1687 965 1717 982
rect 1687 948 1694 965
rect 1711 948 1717 965
rect 1687 931 1717 948
rect 1687 914 1694 931
rect 1711 914 1717 931
rect 1687 897 1717 914
rect 1687 880 1694 897
rect 1711 880 1717 897
rect 1687 863 1717 880
rect 1687 846 1694 863
rect 1711 846 1717 863
rect 1687 829 1717 846
rect 1687 812 1694 829
rect 1711 812 1717 829
rect 1687 795 1717 812
rect 1687 778 1694 795
rect 1711 778 1717 795
rect 1687 761 1717 778
rect 1687 744 1694 761
rect 1711 744 1717 761
rect 1687 727 1717 744
rect 1687 710 1694 727
rect 1711 710 1717 727
rect 1687 693 1717 710
rect 1687 676 1694 693
rect 1711 676 1717 693
rect 1687 659 1717 676
rect 1687 642 1694 659
rect 1711 642 1717 659
rect 1687 625 1717 642
rect 1687 608 1694 625
rect 1711 608 1717 625
rect 1687 591 1717 608
rect 1687 574 1694 591
rect 1711 574 1717 591
rect 1687 557 1717 574
rect 1687 540 1694 557
rect 1711 540 1717 557
rect 1687 523 1717 540
rect 1687 506 1694 523
rect 1711 506 1717 523
rect 1687 489 1717 506
rect 1687 472 1694 489
rect 1711 472 1717 489
rect 1687 455 1717 472
rect 1687 438 1694 455
rect 1711 438 1717 455
rect 1687 421 1717 438
rect 1687 404 1694 421
rect 1711 404 1717 421
rect 1687 387 1717 404
rect 1687 370 1694 387
rect 1711 370 1717 387
rect 1687 353 1717 370
rect 1687 336 1694 353
rect 1711 336 1717 353
rect 1687 319 1717 336
rect 1687 302 1694 319
rect 1711 302 1717 319
rect 1687 285 1717 302
rect 1687 268 1694 285
rect 1711 268 1717 285
rect 1687 251 1717 268
rect 1687 234 1694 251
rect 1711 234 1717 251
rect 1687 217 1717 234
rect 1687 200 1694 217
rect 1711 200 1717 217
rect 1687 183 1717 200
rect 1687 166 1694 183
rect 1711 166 1717 183
rect 1687 150 1717 166
rect 1732 1135 1763 1150
rect 1732 1118 1739 1135
rect 1756 1118 1763 1135
rect 1732 1101 1763 1118
rect 1732 1084 1739 1101
rect 1756 1084 1763 1101
rect 1732 1067 1763 1084
rect 1732 1050 1739 1067
rect 1756 1050 1763 1067
rect 1732 1033 1763 1050
rect 1732 1016 1739 1033
rect 1756 1016 1763 1033
rect 1732 999 1763 1016
rect 1732 982 1740 999
rect 1757 982 1763 999
rect 1732 965 1763 982
rect 1732 948 1740 965
rect 1757 948 1763 965
rect 1732 931 1763 948
rect 1732 914 1740 931
rect 1757 914 1763 931
rect 1732 897 1763 914
rect 1732 880 1740 897
rect 1757 880 1763 897
rect 1732 863 1763 880
rect 1732 846 1740 863
rect 1757 846 1763 863
rect 1732 829 1763 846
rect 1732 812 1740 829
rect 1757 812 1763 829
rect 1732 795 1763 812
rect 1732 778 1740 795
rect 1757 778 1763 795
rect 1732 761 1763 778
rect 1732 744 1740 761
rect 1757 744 1763 761
rect 1732 727 1763 744
rect 1732 710 1740 727
rect 1757 710 1763 727
rect 1732 693 1763 710
rect 1732 676 1740 693
rect 1757 676 1763 693
rect 1732 659 1763 676
rect 1732 642 1740 659
rect 1757 642 1763 659
rect 1732 625 1763 642
rect 1732 608 1740 625
rect 1757 608 1763 625
rect 1732 591 1763 608
rect 1732 574 1740 591
rect 1757 574 1763 591
rect 1732 557 1763 574
rect 1732 540 1740 557
rect 1757 540 1763 557
rect 1732 523 1763 540
rect 1732 506 1740 523
rect 1757 506 1763 523
rect 1732 489 1763 506
rect 1732 472 1740 489
rect 1757 472 1763 489
rect 1732 455 1763 472
rect 1732 438 1740 455
rect 1757 438 1763 455
rect 1732 421 1763 438
rect 1732 404 1740 421
rect 1757 404 1763 421
rect 1732 387 1763 404
rect 1732 370 1740 387
rect 1757 370 1763 387
rect 1732 353 1763 370
rect 1732 336 1740 353
rect 1757 336 1763 353
rect 1732 319 1763 336
rect 1732 302 1740 319
rect 1757 302 1763 319
rect 1732 285 1763 302
rect 1732 268 1740 285
rect 1757 268 1763 285
rect 1732 251 1763 268
rect 1732 234 1740 251
rect 1757 234 1763 251
rect 1732 217 1763 234
rect 1732 200 1740 217
rect 1757 200 1763 217
rect 1732 183 1763 200
rect 1732 166 1740 183
rect 1757 166 1763 183
rect 1732 150 1763 166
rect 1778 1137 1807 1150
rect 1778 1120 1784 1137
rect 1801 1120 1807 1137
rect 1778 1103 1807 1120
rect 1778 1086 1784 1103
rect 1801 1086 1807 1103
rect 1778 1069 1807 1086
rect 1778 1052 1784 1069
rect 1801 1052 1807 1069
rect 1778 1035 1807 1052
rect 1778 1018 1784 1035
rect 1801 1018 1807 1035
rect 1778 1001 1807 1018
rect 1778 984 1784 1001
rect 1801 984 1807 1001
rect 1778 967 1807 984
rect 1778 950 1784 967
rect 1801 950 1807 967
rect 1778 933 1807 950
rect 1778 916 1784 933
rect 1801 916 1807 933
rect 1778 899 1807 916
rect 1778 882 1784 899
rect 1801 882 1807 899
rect 1778 865 1807 882
rect 1778 848 1784 865
rect 1801 848 1807 865
rect 1778 831 1807 848
rect 1778 814 1784 831
rect 1801 814 1807 831
rect 1778 797 1807 814
rect 1778 780 1784 797
rect 1801 780 1807 797
rect 1778 763 1807 780
rect 1778 746 1784 763
rect 1801 746 1807 763
rect 1778 729 1807 746
rect 1778 712 1784 729
rect 1801 712 1807 729
rect 1778 695 1807 712
rect 1778 678 1784 695
rect 1801 678 1807 695
rect 1778 661 1807 678
rect 1778 644 1784 661
rect 1801 644 1807 661
rect 1778 627 1807 644
rect 1778 610 1784 627
rect 1801 610 1807 627
rect 1778 593 1807 610
rect 1778 576 1784 593
rect 1801 576 1807 593
rect 1778 559 1807 576
rect 1778 542 1784 559
rect 1801 542 1807 559
rect 1778 525 1807 542
rect 1778 508 1784 525
rect 1801 508 1807 525
rect 1778 491 1807 508
rect 1778 474 1784 491
rect 1801 474 1807 491
rect 1778 457 1807 474
rect 1778 440 1784 457
rect 1801 440 1807 457
rect 1778 423 1807 440
rect 1778 406 1784 423
rect 1801 406 1807 423
rect 1778 389 1807 406
rect 1778 372 1784 389
rect 1801 372 1807 389
rect 1778 355 1807 372
rect 1778 338 1784 355
rect 1801 338 1807 355
rect 1778 321 1807 338
rect 1778 304 1784 321
rect 1801 304 1807 321
rect 1778 287 1807 304
rect 1778 270 1784 287
rect 1801 270 1807 287
rect 1778 253 1807 270
rect 1778 236 1784 253
rect 1801 236 1807 253
rect 1778 219 1807 236
rect 1778 202 1784 219
rect 1801 202 1807 219
rect 1778 185 1807 202
rect 1778 168 1784 185
rect 1801 168 1807 185
rect 1778 150 1807 168
rect 1822 1135 1852 1150
rect 1822 1118 1828 1135
rect 1845 1118 1852 1135
rect 1822 1101 1852 1118
rect 1822 1084 1828 1101
rect 1845 1084 1852 1101
rect 1822 1067 1852 1084
rect 1822 1050 1828 1067
rect 1845 1050 1852 1067
rect 1822 1033 1852 1050
rect 1822 1016 1828 1033
rect 1845 1016 1852 1033
rect 1822 999 1852 1016
rect 1822 982 1829 999
rect 1846 982 1852 999
rect 1822 965 1852 982
rect 1822 948 1829 965
rect 1846 948 1852 965
rect 1822 931 1852 948
rect 1822 914 1829 931
rect 1846 914 1852 931
rect 1822 897 1852 914
rect 1822 880 1829 897
rect 1846 880 1852 897
rect 1822 863 1852 880
rect 1822 846 1829 863
rect 1846 846 1852 863
rect 1822 829 1852 846
rect 1822 812 1829 829
rect 1846 812 1852 829
rect 1822 795 1852 812
rect 1822 778 1829 795
rect 1846 778 1852 795
rect 1822 761 1852 778
rect 1822 744 1829 761
rect 1846 744 1852 761
rect 1822 727 1852 744
rect 1822 710 1829 727
rect 1846 710 1852 727
rect 1822 693 1852 710
rect 1822 676 1829 693
rect 1846 676 1852 693
rect 1822 659 1852 676
rect 1822 642 1829 659
rect 1846 642 1852 659
rect 1822 625 1852 642
rect 1822 608 1829 625
rect 1846 608 1852 625
rect 1822 591 1852 608
rect 1822 574 1829 591
rect 1846 574 1852 591
rect 1822 557 1852 574
rect 1822 540 1829 557
rect 1846 540 1852 557
rect 1822 523 1852 540
rect 1822 506 1829 523
rect 1846 506 1852 523
rect 1822 489 1852 506
rect 1822 472 1829 489
rect 1846 472 1852 489
rect 1822 455 1852 472
rect 1822 438 1829 455
rect 1846 438 1852 455
rect 1822 421 1852 438
rect 1822 404 1829 421
rect 1846 404 1852 421
rect 1822 387 1852 404
rect 1822 370 1829 387
rect 1846 370 1852 387
rect 1822 353 1852 370
rect 1822 336 1829 353
rect 1846 336 1852 353
rect 1822 319 1852 336
rect 1822 302 1829 319
rect 1846 302 1852 319
rect 1822 285 1852 302
rect 1822 268 1829 285
rect 1846 268 1852 285
rect 1822 251 1852 268
rect 1822 234 1829 251
rect 1846 234 1852 251
rect 1822 217 1852 234
rect 1822 200 1829 217
rect 1846 200 1852 217
rect 1822 183 1852 200
rect 1822 166 1829 183
rect 1846 166 1852 183
rect 1822 150 1852 166
rect 1867 1135 1897 1150
rect 1867 1118 1873 1135
rect 1890 1118 1897 1135
rect 1867 1101 1897 1118
rect 1867 1084 1873 1101
rect 1890 1084 1897 1101
rect 1867 1067 1897 1084
rect 1867 1050 1873 1067
rect 1890 1050 1897 1067
rect 1867 1033 1897 1050
rect 1867 1016 1873 1033
rect 1890 1016 1897 1033
rect 1867 999 1897 1016
rect 1867 982 1874 999
rect 1891 982 1897 999
rect 1867 965 1897 982
rect 1867 948 1874 965
rect 1891 948 1897 965
rect 1867 931 1897 948
rect 1867 914 1874 931
rect 1891 914 1897 931
rect 1867 897 1897 914
rect 1867 880 1874 897
rect 1891 880 1897 897
rect 1867 863 1897 880
rect 1867 846 1874 863
rect 1891 846 1897 863
rect 1867 829 1897 846
rect 1867 812 1874 829
rect 1891 812 1897 829
rect 1867 795 1897 812
rect 1867 778 1874 795
rect 1891 778 1897 795
rect 1867 761 1897 778
rect 1867 744 1874 761
rect 1891 744 1897 761
rect 1867 727 1897 744
rect 1867 710 1874 727
rect 1891 710 1897 727
rect 1867 693 1897 710
rect 1867 676 1874 693
rect 1891 676 1897 693
rect 1867 659 1897 676
rect 1867 642 1874 659
rect 1891 642 1897 659
rect 1867 625 1897 642
rect 1867 608 1874 625
rect 1891 608 1897 625
rect 1867 591 1897 608
rect 1867 574 1874 591
rect 1891 574 1897 591
rect 1867 557 1897 574
rect 1867 540 1874 557
rect 1891 540 1897 557
rect 1867 523 1897 540
rect 1867 506 1874 523
rect 1891 506 1897 523
rect 1867 489 1897 506
rect 1867 472 1874 489
rect 1891 472 1897 489
rect 1867 455 1897 472
rect 1867 438 1874 455
rect 1891 438 1897 455
rect 1867 421 1897 438
rect 1867 404 1874 421
rect 1891 404 1897 421
rect 1867 387 1897 404
rect 1867 370 1874 387
rect 1891 370 1897 387
rect 1867 353 1897 370
rect 1867 336 1874 353
rect 1891 336 1897 353
rect 1867 319 1897 336
rect 1867 302 1874 319
rect 1891 302 1897 319
rect 1867 285 1897 302
rect 1867 268 1874 285
rect 1891 268 1897 285
rect 1867 251 1897 268
rect 1867 234 1874 251
rect 1891 234 1897 251
rect 1867 217 1897 234
rect 1867 200 1874 217
rect 1891 200 1897 217
rect 1867 183 1897 200
rect 1867 166 1874 183
rect 1891 166 1897 183
rect 1867 150 1897 166
rect 1912 1135 1942 1150
rect 1912 1118 1918 1135
rect 1935 1118 1942 1135
rect 1912 1101 1942 1118
rect 1912 1084 1918 1101
rect 1935 1084 1942 1101
rect 1912 1067 1942 1084
rect 1912 1050 1918 1067
rect 1935 1050 1942 1067
rect 1912 1033 1942 1050
rect 1912 1016 1918 1033
rect 1935 1016 1942 1033
rect 1912 999 1942 1016
rect 1912 982 1919 999
rect 1936 982 1942 999
rect 1912 965 1942 982
rect 1912 948 1919 965
rect 1936 948 1942 965
rect 1912 931 1942 948
rect 1912 914 1919 931
rect 1936 914 1942 931
rect 1912 897 1942 914
rect 1912 880 1919 897
rect 1936 880 1942 897
rect 1912 863 1942 880
rect 1912 846 1919 863
rect 1936 846 1942 863
rect 1912 829 1942 846
rect 1912 812 1919 829
rect 1936 812 1942 829
rect 1912 795 1942 812
rect 1912 778 1919 795
rect 1936 778 1942 795
rect 1912 761 1942 778
rect 1912 744 1919 761
rect 1936 744 1942 761
rect 1912 727 1942 744
rect 1912 710 1919 727
rect 1936 710 1942 727
rect 1912 693 1942 710
rect 1912 676 1919 693
rect 1936 676 1942 693
rect 1912 659 1942 676
rect 1912 642 1919 659
rect 1936 642 1942 659
rect 1912 625 1942 642
rect 1912 608 1919 625
rect 1936 608 1942 625
rect 1912 591 1942 608
rect 1912 574 1919 591
rect 1936 574 1942 591
rect 1912 557 1942 574
rect 1912 540 1919 557
rect 1936 540 1942 557
rect 1912 523 1942 540
rect 1912 506 1919 523
rect 1936 506 1942 523
rect 1912 489 1942 506
rect 1912 472 1919 489
rect 1936 472 1942 489
rect 1912 455 1942 472
rect 1912 438 1919 455
rect 1936 438 1942 455
rect 1912 421 1942 438
rect 1912 404 1919 421
rect 1936 404 1942 421
rect 1912 387 1942 404
rect 1912 370 1919 387
rect 1936 370 1942 387
rect 1912 353 1942 370
rect 1912 336 1919 353
rect 1936 336 1942 353
rect 1912 319 1942 336
rect 1912 302 1919 319
rect 1936 302 1942 319
rect 1912 285 1942 302
rect 1912 268 1919 285
rect 1936 268 1942 285
rect 1912 251 1942 268
rect 1912 234 1919 251
rect 1936 234 1942 251
rect 1912 217 1942 234
rect 1912 200 1919 217
rect 1936 200 1942 217
rect 1912 183 1942 200
rect 1912 166 1919 183
rect 1936 166 1942 183
rect 1912 150 1942 166
rect 1957 1135 1987 1150
rect 1957 1118 1963 1135
rect 1980 1118 1987 1135
rect 1957 1101 1987 1118
rect 1957 1084 1963 1101
rect 1980 1084 1987 1101
rect 1957 1067 1987 1084
rect 1957 1050 1963 1067
rect 1980 1050 1987 1067
rect 1957 1033 1987 1050
rect 1957 1016 1963 1033
rect 1980 1016 1987 1033
rect 1957 999 1987 1016
rect 1957 982 1964 999
rect 1981 982 1987 999
rect 1957 965 1987 982
rect 1957 948 1964 965
rect 1981 948 1987 965
rect 1957 931 1987 948
rect 1957 914 1964 931
rect 1981 914 1987 931
rect 1957 897 1987 914
rect 1957 880 1964 897
rect 1981 880 1987 897
rect 1957 863 1987 880
rect 1957 846 1964 863
rect 1981 846 1987 863
rect 1957 829 1987 846
rect 1957 812 1964 829
rect 1981 812 1987 829
rect 1957 795 1987 812
rect 1957 778 1964 795
rect 1981 778 1987 795
rect 1957 761 1987 778
rect 1957 744 1964 761
rect 1981 744 1987 761
rect 1957 727 1987 744
rect 1957 710 1964 727
rect 1981 710 1987 727
rect 1957 693 1987 710
rect 1957 676 1964 693
rect 1981 676 1987 693
rect 1957 659 1987 676
rect 1957 642 1964 659
rect 1981 642 1987 659
rect 1957 625 1987 642
rect 1957 608 1964 625
rect 1981 608 1987 625
rect 1957 591 1987 608
rect 1957 574 1964 591
rect 1981 574 1987 591
rect 1957 557 1987 574
rect 1957 540 1964 557
rect 1981 540 1987 557
rect 1957 523 1987 540
rect 1957 506 1964 523
rect 1981 506 1987 523
rect 1957 489 1987 506
rect 1957 472 1964 489
rect 1981 472 1987 489
rect 1957 455 1987 472
rect 1957 438 1964 455
rect 1981 438 1987 455
rect 1957 421 1987 438
rect 1957 404 1964 421
rect 1981 404 1987 421
rect 1957 387 1987 404
rect 1957 370 1964 387
rect 1981 370 1987 387
rect 1957 353 1987 370
rect 1957 336 1964 353
rect 1981 336 1987 353
rect 1957 319 1987 336
rect 1957 302 1964 319
rect 1981 302 1987 319
rect 1957 285 1987 302
rect 1957 268 1964 285
rect 1981 268 1987 285
rect 1957 251 1987 268
rect 1957 234 1964 251
rect 1981 234 1987 251
rect 1957 217 1987 234
rect 1957 200 1964 217
rect 1981 200 1987 217
rect 1957 183 1987 200
rect 1957 166 1964 183
rect 1981 166 1987 183
rect 1957 150 1987 166
rect 2002 1135 2032 1150
rect 2002 1118 2008 1135
rect 2025 1118 2032 1135
rect 2002 1101 2032 1118
rect 2002 1084 2008 1101
rect 2025 1084 2032 1101
rect 2002 1067 2032 1084
rect 2002 1050 2008 1067
rect 2025 1050 2032 1067
rect 2002 1033 2032 1050
rect 2002 1016 2008 1033
rect 2025 1016 2032 1033
rect 2002 999 2032 1016
rect 2002 982 2009 999
rect 2026 982 2032 999
rect 2002 965 2032 982
rect 2002 948 2009 965
rect 2026 948 2032 965
rect 2002 931 2032 948
rect 2002 914 2009 931
rect 2026 914 2032 931
rect 2002 897 2032 914
rect 2002 880 2009 897
rect 2026 880 2032 897
rect 2002 863 2032 880
rect 2002 846 2009 863
rect 2026 846 2032 863
rect 2002 829 2032 846
rect 2002 812 2009 829
rect 2026 812 2032 829
rect 2002 795 2032 812
rect 2002 778 2009 795
rect 2026 778 2032 795
rect 2002 761 2032 778
rect 2002 744 2009 761
rect 2026 744 2032 761
rect 2002 727 2032 744
rect 2002 710 2009 727
rect 2026 710 2032 727
rect 2002 693 2032 710
rect 2002 676 2009 693
rect 2026 676 2032 693
rect 2002 659 2032 676
rect 2002 642 2009 659
rect 2026 642 2032 659
rect 2002 625 2032 642
rect 2002 608 2009 625
rect 2026 608 2032 625
rect 2002 591 2032 608
rect 2002 574 2009 591
rect 2026 574 2032 591
rect 2002 557 2032 574
rect 2002 540 2009 557
rect 2026 540 2032 557
rect 2002 523 2032 540
rect 2002 506 2009 523
rect 2026 506 2032 523
rect 2002 489 2032 506
rect 2002 472 2009 489
rect 2026 472 2032 489
rect 2002 455 2032 472
rect 2002 438 2009 455
rect 2026 438 2032 455
rect 2002 421 2032 438
rect 2002 404 2009 421
rect 2026 404 2032 421
rect 2002 387 2032 404
rect 2002 370 2009 387
rect 2026 370 2032 387
rect 2002 353 2032 370
rect 2002 336 2009 353
rect 2026 336 2032 353
rect 2002 319 2032 336
rect 2002 302 2009 319
rect 2026 302 2032 319
rect 2002 285 2032 302
rect 2002 268 2009 285
rect 2026 268 2032 285
rect 2002 251 2032 268
rect 2002 234 2009 251
rect 2026 234 2032 251
rect 2002 217 2032 234
rect 2002 200 2009 217
rect 2026 200 2032 217
rect 2002 183 2032 200
rect 2002 166 2009 183
rect 2026 166 2032 183
rect 2002 150 2032 166
rect 2047 1135 2077 1150
rect 2047 1118 2053 1135
rect 2070 1118 2077 1135
rect 2047 1101 2077 1118
rect 2047 1084 2053 1101
rect 2070 1084 2077 1101
rect 2047 1067 2077 1084
rect 2047 1050 2053 1067
rect 2070 1050 2077 1067
rect 2047 1033 2077 1050
rect 2047 1016 2053 1033
rect 2070 1016 2077 1033
rect 2047 999 2077 1016
rect 2047 982 2054 999
rect 2071 982 2077 999
rect 2047 965 2077 982
rect 2047 948 2054 965
rect 2071 948 2077 965
rect 2047 931 2077 948
rect 2047 914 2054 931
rect 2071 914 2077 931
rect 2047 897 2077 914
rect 2047 880 2054 897
rect 2071 880 2077 897
rect 2047 863 2077 880
rect 2047 846 2054 863
rect 2071 846 2077 863
rect 2047 829 2077 846
rect 2047 812 2054 829
rect 2071 812 2077 829
rect 2047 795 2077 812
rect 2047 778 2054 795
rect 2071 778 2077 795
rect 2047 761 2077 778
rect 2047 744 2054 761
rect 2071 744 2077 761
rect 2047 727 2077 744
rect 2047 710 2054 727
rect 2071 710 2077 727
rect 2047 693 2077 710
rect 2047 676 2054 693
rect 2071 676 2077 693
rect 2047 659 2077 676
rect 2047 642 2054 659
rect 2071 642 2077 659
rect 2047 625 2077 642
rect 2047 608 2054 625
rect 2071 608 2077 625
rect 2047 591 2077 608
rect 2047 574 2054 591
rect 2071 574 2077 591
rect 2047 557 2077 574
rect 2047 540 2054 557
rect 2071 540 2077 557
rect 2047 523 2077 540
rect 2047 506 2054 523
rect 2071 506 2077 523
rect 2047 489 2077 506
rect 2047 472 2054 489
rect 2071 472 2077 489
rect 2047 455 2077 472
rect 2047 438 2054 455
rect 2071 438 2077 455
rect 2047 421 2077 438
rect 2047 404 2054 421
rect 2071 404 2077 421
rect 2047 387 2077 404
rect 2047 370 2054 387
rect 2071 370 2077 387
rect 2047 353 2077 370
rect 2047 336 2054 353
rect 2071 336 2077 353
rect 2047 319 2077 336
rect 2047 302 2054 319
rect 2071 302 2077 319
rect 2047 285 2077 302
rect 2047 268 2054 285
rect 2071 268 2077 285
rect 2047 251 2077 268
rect 2047 234 2054 251
rect 2071 234 2077 251
rect 2047 217 2077 234
rect 2047 200 2054 217
rect 2071 200 2077 217
rect 2047 183 2077 200
rect 2047 166 2054 183
rect 2071 166 2077 183
rect 2047 150 2077 166
rect 2092 1135 2122 1150
rect 2092 1118 2098 1135
rect 2115 1118 2122 1135
rect 2092 1101 2122 1118
rect 2092 1084 2098 1101
rect 2115 1084 2122 1101
rect 2092 1067 2122 1084
rect 2092 1050 2098 1067
rect 2115 1050 2122 1067
rect 2092 1033 2122 1050
rect 2092 1016 2098 1033
rect 2115 1016 2122 1033
rect 2092 999 2122 1016
rect 2092 982 2099 999
rect 2116 982 2122 999
rect 2092 965 2122 982
rect 2092 948 2099 965
rect 2116 948 2122 965
rect 2092 931 2122 948
rect 2092 914 2099 931
rect 2116 914 2122 931
rect 2092 897 2122 914
rect 2092 880 2099 897
rect 2116 880 2122 897
rect 2092 863 2122 880
rect 2092 846 2099 863
rect 2116 846 2122 863
rect 2092 829 2122 846
rect 2092 812 2099 829
rect 2116 812 2122 829
rect 2092 795 2122 812
rect 2092 778 2099 795
rect 2116 778 2122 795
rect 2092 761 2122 778
rect 2092 744 2099 761
rect 2116 744 2122 761
rect 2092 727 2122 744
rect 2092 710 2099 727
rect 2116 710 2122 727
rect 2092 693 2122 710
rect 2092 676 2099 693
rect 2116 676 2122 693
rect 2092 659 2122 676
rect 2092 642 2099 659
rect 2116 642 2122 659
rect 2092 625 2122 642
rect 2092 608 2099 625
rect 2116 608 2122 625
rect 2092 591 2122 608
rect 2092 574 2099 591
rect 2116 574 2122 591
rect 2092 557 2122 574
rect 2092 540 2099 557
rect 2116 540 2122 557
rect 2092 523 2122 540
rect 2092 506 2099 523
rect 2116 506 2122 523
rect 2092 489 2122 506
rect 2092 472 2099 489
rect 2116 472 2122 489
rect 2092 455 2122 472
rect 2092 438 2099 455
rect 2116 438 2122 455
rect 2092 421 2122 438
rect 2092 404 2099 421
rect 2116 404 2122 421
rect 2092 387 2122 404
rect 2092 370 2099 387
rect 2116 370 2122 387
rect 2092 353 2122 370
rect 2092 336 2099 353
rect 2116 336 2122 353
rect 2092 319 2122 336
rect 2092 302 2099 319
rect 2116 302 2122 319
rect 2092 285 2122 302
rect 2092 268 2099 285
rect 2116 268 2122 285
rect 2092 251 2122 268
rect 2092 234 2099 251
rect 2116 234 2122 251
rect 2092 217 2122 234
rect 2092 200 2099 217
rect 2116 200 2122 217
rect 2092 183 2122 200
rect 2092 166 2099 183
rect 2116 166 2122 183
rect 2092 150 2122 166
rect 2137 1137 2166 1150
rect 2137 1120 2143 1137
rect 2160 1120 2166 1137
rect 2137 1103 2166 1120
rect 2137 1086 2143 1103
rect 2160 1086 2166 1103
rect 2137 1069 2166 1086
rect 2137 1052 2143 1069
rect 2160 1052 2166 1069
rect 2137 1035 2166 1052
rect 2137 1018 2143 1035
rect 2160 1018 2166 1035
rect 2137 1001 2166 1018
rect 2137 984 2143 1001
rect 2160 984 2166 1001
rect 2137 967 2166 984
rect 2137 950 2143 967
rect 2160 950 2166 967
rect 2137 933 2166 950
rect 2137 916 2143 933
rect 2160 916 2166 933
rect 2137 899 2166 916
rect 2137 882 2143 899
rect 2160 882 2166 899
rect 2137 865 2166 882
rect 2137 848 2143 865
rect 2160 848 2166 865
rect 2137 831 2166 848
rect 2137 814 2143 831
rect 2160 814 2166 831
rect 2137 797 2166 814
rect 2137 780 2143 797
rect 2160 780 2166 797
rect 2137 763 2166 780
rect 2137 746 2143 763
rect 2160 746 2166 763
rect 2137 729 2166 746
rect 2137 712 2143 729
rect 2160 712 2166 729
rect 2137 695 2166 712
rect 2137 678 2143 695
rect 2160 678 2166 695
rect 2137 661 2166 678
rect 2137 644 2143 661
rect 2160 644 2166 661
rect 2137 627 2166 644
rect 2137 610 2143 627
rect 2160 610 2166 627
rect 2137 593 2166 610
rect 2137 576 2143 593
rect 2160 576 2166 593
rect 2137 559 2166 576
rect 2137 542 2143 559
rect 2160 542 2166 559
rect 2137 525 2166 542
rect 2137 508 2143 525
rect 2160 508 2166 525
rect 2137 491 2166 508
rect 2137 474 2143 491
rect 2160 474 2166 491
rect 2137 457 2166 474
rect 2137 440 2143 457
rect 2160 440 2166 457
rect 2137 423 2166 440
rect 2137 406 2143 423
rect 2160 406 2166 423
rect 2137 389 2166 406
rect 2137 372 2143 389
rect 2160 372 2166 389
rect 2137 355 2166 372
rect 2137 338 2143 355
rect 2160 338 2166 355
rect 2137 321 2166 338
rect 2137 304 2143 321
rect 2160 304 2166 321
rect 2137 287 2166 304
rect 2137 270 2143 287
rect 2160 270 2166 287
rect 2137 253 2166 270
rect 2137 236 2143 253
rect 2160 236 2166 253
rect 2137 219 2166 236
rect 2137 202 2143 219
rect 2160 202 2166 219
rect 2137 185 2166 202
rect 2137 168 2143 185
rect 2160 168 2166 185
rect 2137 150 2166 168
rect 2181 1135 2211 1150
rect 2181 1118 2187 1135
rect 2204 1118 2211 1135
rect 2181 1101 2211 1118
rect 2181 1084 2187 1101
rect 2204 1084 2211 1101
rect 2181 1067 2211 1084
rect 2181 1050 2187 1067
rect 2204 1050 2211 1067
rect 2181 1033 2211 1050
rect 2181 1016 2187 1033
rect 2204 1016 2211 1033
rect 2181 999 2211 1016
rect 2181 982 2188 999
rect 2205 982 2211 999
rect 2181 965 2211 982
rect 2181 948 2188 965
rect 2205 948 2211 965
rect 2181 931 2211 948
rect 2181 914 2188 931
rect 2205 914 2211 931
rect 2181 897 2211 914
rect 2181 880 2188 897
rect 2205 880 2211 897
rect 2181 863 2211 880
rect 2181 846 2188 863
rect 2205 846 2211 863
rect 2181 829 2211 846
rect 2181 812 2188 829
rect 2205 812 2211 829
rect 2181 795 2211 812
rect 2181 778 2188 795
rect 2205 778 2211 795
rect 2181 761 2211 778
rect 2181 744 2188 761
rect 2205 744 2211 761
rect 2181 727 2211 744
rect 2181 710 2188 727
rect 2205 710 2211 727
rect 2181 693 2211 710
rect 2181 676 2188 693
rect 2205 676 2211 693
rect 2181 659 2211 676
rect 2181 642 2188 659
rect 2205 642 2211 659
rect 2181 625 2211 642
rect 2181 608 2188 625
rect 2205 608 2211 625
rect 2181 591 2211 608
rect 2181 574 2188 591
rect 2205 574 2211 591
rect 2181 557 2211 574
rect 2181 540 2188 557
rect 2205 540 2211 557
rect 2181 523 2211 540
rect 2181 506 2188 523
rect 2205 506 2211 523
rect 2181 489 2211 506
rect 2181 472 2188 489
rect 2205 472 2211 489
rect 2181 455 2211 472
rect 2181 438 2188 455
rect 2205 438 2211 455
rect 2181 421 2211 438
rect 2181 404 2188 421
rect 2205 404 2211 421
rect 2181 387 2211 404
rect 2181 370 2188 387
rect 2205 370 2211 387
rect 2181 353 2211 370
rect 2181 336 2188 353
rect 2205 336 2211 353
rect 2181 319 2211 336
rect 2181 302 2188 319
rect 2205 302 2211 319
rect 2181 285 2211 302
rect 2181 268 2188 285
rect 2205 268 2211 285
rect 2181 251 2211 268
rect 2181 234 2188 251
rect 2205 234 2211 251
rect 2181 217 2211 234
rect 2181 200 2188 217
rect 2205 200 2211 217
rect 2181 183 2211 200
rect 2181 166 2188 183
rect 2205 166 2211 183
rect 2181 150 2211 166
rect 2226 1135 2256 1150
rect 2226 1118 2232 1135
rect 2249 1118 2256 1135
rect 2226 1101 2256 1118
rect 2226 1084 2232 1101
rect 2249 1084 2256 1101
rect 2226 1067 2256 1084
rect 2226 1050 2232 1067
rect 2249 1050 2256 1067
rect 2226 1033 2256 1050
rect 2226 1016 2232 1033
rect 2249 1016 2256 1033
rect 2226 999 2256 1016
rect 2226 982 2233 999
rect 2250 982 2256 999
rect 2226 965 2256 982
rect 2226 948 2233 965
rect 2250 948 2256 965
rect 2226 931 2256 948
rect 2226 914 2233 931
rect 2250 914 2256 931
rect 2226 897 2256 914
rect 2226 880 2233 897
rect 2250 880 2256 897
rect 2226 863 2256 880
rect 2226 846 2233 863
rect 2250 846 2256 863
rect 2226 829 2256 846
rect 2226 812 2233 829
rect 2250 812 2256 829
rect 2226 795 2256 812
rect 2226 778 2233 795
rect 2250 778 2256 795
rect 2226 761 2256 778
rect 2226 744 2233 761
rect 2250 744 2256 761
rect 2226 727 2256 744
rect 2226 710 2233 727
rect 2250 710 2256 727
rect 2226 693 2256 710
rect 2226 676 2233 693
rect 2250 676 2256 693
rect 2226 659 2256 676
rect 2226 642 2233 659
rect 2250 642 2256 659
rect 2226 625 2256 642
rect 2226 608 2233 625
rect 2250 608 2256 625
rect 2226 591 2256 608
rect 2226 574 2233 591
rect 2250 574 2256 591
rect 2226 557 2256 574
rect 2226 540 2233 557
rect 2250 540 2256 557
rect 2226 523 2256 540
rect 2226 506 2233 523
rect 2250 506 2256 523
rect 2226 489 2256 506
rect 2226 472 2233 489
rect 2250 472 2256 489
rect 2226 455 2256 472
rect 2226 438 2233 455
rect 2250 438 2256 455
rect 2226 421 2256 438
rect 2226 404 2233 421
rect 2250 404 2256 421
rect 2226 387 2256 404
rect 2226 370 2233 387
rect 2250 370 2256 387
rect 2226 353 2256 370
rect 2226 336 2233 353
rect 2250 336 2256 353
rect 2226 319 2256 336
rect 2226 302 2233 319
rect 2250 302 2256 319
rect 2226 285 2256 302
rect 2226 268 2233 285
rect 2250 268 2256 285
rect 2226 251 2256 268
rect 2226 234 2233 251
rect 2250 234 2256 251
rect 2226 217 2256 234
rect 2226 200 2233 217
rect 2250 200 2256 217
rect 2226 183 2256 200
rect 2226 166 2233 183
rect 2250 166 2256 183
rect 2226 150 2256 166
rect 2271 1135 2301 1150
rect 2271 1118 2277 1135
rect 2294 1118 2301 1135
rect 2271 1101 2301 1118
rect 2271 1084 2277 1101
rect 2294 1084 2301 1101
rect 2271 1067 2301 1084
rect 2271 1050 2277 1067
rect 2294 1050 2301 1067
rect 2271 1033 2301 1050
rect 2271 1016 2277 1033
rect 2294 1016 2301 1033
rect 2271 999 2301 1016
rect 2271 982 2278 999
rect 2295 982 2301 999
rect 2271 965 2301 982
rect 2271 948 2278 965
rect 2295 948 2301 965
rect 2271 931 2301 948
rect 2271 914 2278 931
rect 2295 914 2301 931
rect 2271 897 2301 914
rect 2271 880 2278 897
rect 2295 880 2301 897
rect 2271 863 2301 880
rect 2271 846 2278 863
rect 2295 846 2301 863
rect 2271 829 2301 846
rect 2271 812 2278 829
rect 2295 812 2301 829
rect 2271 795 2301 812
rect 2271 778 2278 795
rect 2295 778 2301 795
rect 2271 761 2301 778
rect 2271 744 2278 761
rect 2295 744 2301 761
rect 2271 727 2301 744
rect 2271 710 2278 727
rect 2295 710 2301 727
rect 2271 693 2301 710
rect 2271 676 2278 693
rect 2295 676 2301 693
rect 2271 659 2301 676
rect 2271 642 2278 659
rect 2295 642 2301 659
rect 2271 625 2301 642
rect 2271 608 2278 625
rect 2295 608 2301 625
rect 2271 591 2301 608
rect 2271 574 2278 591
rect 2295 574 2301 591
rect 2271 557 2301 574
rect 2271 540 2278 557
rect 2295 540 2301 557
rect 2271 523 2301 540
rect 2271 506 2278 523
rect 2295 506 2301 523
rect 2271 489 2301 506
rect 2271 472 2278 489
rect 2295 472 2301 489
rect 2271 455 2301 472
rect 2271 438 2278 455
rect 2295 438 2301 455
rect 2271 421 2301 438
rect 2271 404 2278 421
rect 2295 404 2301 421
rect 2271 387 2301 404
rect 2271 370 2278 387
rect 2295 370 2301 387
rect 2271 353 2301 370
rect 2271 336 2278 353
rect 2295 336 2301 353
rect 2271 319 2301 336
rect 2271 302 2278 319
rect 2295 302 2301 319
rect 2271 285 2301 302
rect 2271 268 2278 285
rect 2295 268 2301 285
rect 2271 251 2301 268
rect 2271 234 2278 251
rect 2295 234 2301 251
rect 2271 217 2301 234
rect 2271 200 2278 217
rect 2295 200 2301 217
rect 2271 183 2301 200
rect 2271 166 2278 183
rect 2295 166 2301 183
rect 2271 150 2301 166
rect 2316 1135 2346 1150
rect 2316 1118 2322 1135
rect 2339 1118 2346 1135
rect 2316 1101 2346 1118
rect 2316 1084 2322 1101
rect 2339 1084 2346 1101
rect 2316 1067 2346 1084
rect 2316 1050 2322 1067
rect 2339 1050 2346 1067
rect 2316 1033 2346 1050
rect 2316 1016 2322 1033
rect 2339 1016 2346 1033
rect 2316 999 2346 1016
rect 2316 982 2323 999
rect 2340 982 2346 999
rect 2316 965 2346 982
rect 2316 948 2323 965
rect 2340 948 2346 965
rect 2316 931 2346 948
rect 2316 914 2323 931
rect 2340 914 2346 931
rect 2316 897 2346 914
rect 2316 880 2323 897
rect 2340 880 2346 897
rect 2316 863 2346 880
rect 2316 846 2323 863
rect 2340 846 2346 863
rect 2316 829 2346 846
rect 2316 812 2323 829
rect 2340 812 2346 829
rect 2316 795 2346 812
rect 2316 778 2323 795
rect 2340 778 2346 795
rect 2316 761 2346 778
rect 2316 744 2323 761
rect 2340 744 2346 761
rect 2316 727 2346 744
rect 2316 710 2323 727
rect 2340 710 2346 727
rect 2316 693 2346 710
rect 2316 676 2323 693
rect 2340 676 2346 693
rect 2316 659 2346 676
rect 2316 642 2323 659
rect 2340 642 2346 659
rect 2316 625 2346 642
rect 2316 608 2323 625
rect 2340 608 2346 625
rect 2316 591 2346 608
rect 2316 574 2323 591
rect 2340 574 2346 591
rect 2316 557 2346 574
rect 2316 540 2323 557
rect 2340 540 2346 557
rect 2316 523 2346 540
rect 2316 506 2323 523
rect 2340 506 2346 523
rect 2316 489 2346 506
rect 2316 472 2323 489
rect 2340 472 2346 489
rect 2316 455 2346 472
rect 2316 438 2323 455
rect 2340 438 2346 455
rect 2316 421 2346 438
rect 2316 404 2323 421
rect 2340 404 2346 421
rect 2316 387 2346 404
rect 2316 370 2323 387
rect 2340 370 2346 387
rect 2316 353 2346 370
rect 2316 336 2323 353
rect 2340 336 2346 353
rect 2316 319 2346 336
rect 2316 302 2323 319
rect 2340 302 2346 319
rect 2316 285 2346 302
rect 2316 268 2323 285
rect 2340 268 2346 285
rect 2316 251 2346 268
rect 2316 234 2323 251
rect 2340 234 2346 251
rect 2316 217 2346 234
rect 2316 200 2323 217
rect 2340 200 2346 217
rect 2316 183 2346 200
rect 2316 166 2323 183
rect 2340 166 2346 183
rect 2316 150 2346 166
rect 2361 1135 2391 1150
rect 2361 1118 2367 1135
rect 2384 1118 2391 1135
rect 2361 1101 2391 1118
rect 2361 1084 2367 1101
rect 2384 1084 2391 1101
rect 2361 1067 2391 1084
rect 2361 1050 2367 1067
rect 2384 1050 2391 1067
rect 2361 1033 2391 1050
rect 2361 1016 2367 1033
rect 2384 1016 2391 1033
rect 2361 999 2391 1016
rect 2361 982 2368 999
rect 2385 982 2391 999
rect 2361 965 2391 982
rect 2361 948 2368 965
rect 2385 948 2391 965
rect 2361 931 2391 948
rect 2361 914 2368 931
rect 2385 914 2391 931
rect 2361 897 2391 914
rect 2361 880 2368 897
rect 2385 880 2391 897
rect 2361 863 2391 880
rect 2361 846 2368 863
rect 2385 846 2391 863
rect 2361 829 2391 846
rect 2361 812 2368 829
rect 2385 812 2391 829
rect 2361 795 2391 812
rect 2361 778 2368 795
rect 2385 778 2391 795
rect 2361 761 2391 778
rect 2361 744 2368 761
rect 2385 744 2391 761
rect 2361 727 2391 744
rect 2361 710 2368 727
rect 2385 710 2391 727
rect 2361 693 2391 710
rect 2361 676 2368 693
rect 2385 676 2391 693
rect 2361 659 2391 676
rect 2361 642 2368 659
rect 2385 642 2391 659
rect 2361 625 2391 642
rect 2361 608 2368 625
rect 2385 608 2391 625
rect 2361 591 2391 608
rect 2361 574 2368 591
rect 2385 574 2391 591
rect 2361 557 2391 574
rect 2361 540 2368 557
rect 2385 540 2391 557
rect 2361 523 2391 540
rect 2361 506 2368 523
rect 2385 506 2391 523
rect 2361 489 2391 506
rect 2361 472 2368 489
rect 2385 472 2391 489
rect 2361 455 2391 472
rect 2361 438 2368 455
rect 2385 438 2391 455
rect 2361 421 2391 438
rect 2361 404 2368 421
rect 2385 404 2391 421
rect 2361 387 2391 404
rect 2361 370 2368 387
rect 2385 370 2391 387
rect 2361 353 2391 370
rect 2361 336 2368 353
rect 2385 336 2391 353
rect 2361 319 2391 336
rect 2361 302 2368 319
rect 2385 302 2391 319
rect 2361 285 2391 302
rect 2361 268 2368 285
rect 2385 268 2391 285
rect 2361 251 2391 268
rect 2361 234 2368 251
rect 2385 234 2391 251
rect 2361 217 2391 234
rect 2361 200 2368 217
rect 2385 200 2391 217
rect 2361 183 2391 200
rect 2361 166 2368 183
rect 2385 166 2391 183
rect 2361 150 2391 166
rect 2406 1135 2436 1150
rect 2406 1118 2412 1135
rect 2429 1118 2436 1135
rect 2406 1101 2436 1118
rect 2406 1084 2412 1101
rect 2429 1084 2436 1101
rect 2406 1067 2436 1084
rect 2406 1050 2412 1067
rect 2429 1050 2436 1067
rect 2406 1033 2436 1050
rect 2406 1016 2412 1033
rect 2429 1016 2436 1033
rect 2406 999 2436 1016
rect 2406 982 2413 999
rect 2430 982 2436 999
rect 2406 965 2436 982
rect 2406 948 2413 965
rect 2430 948 2436 965
rect 2406 931 2436 948
rect 2406 914 2413 931
rect 2430 914 2436 931
rect 2406 897 2436 914
rect 2406 880 2413 897
rect 2430 880 2436 897
rect 2406 863 2436 880
rect 2406 846 2413 863
rect 2430 846 2436 863
rect 2406 829 2436 846
rect 2406 812 2413 829
rect 2430 812 2436 829
rect 2406 795 2436 812
rect 2406 778 2413 795
rect 2430 778 2436 795
rect 2406 761 2436 778
rect 2406 744 2413 761
rect 2430 744 2436 761
rect 2406 727 2436 744
rect 2406 710 2413 727
rect 2430 710 2436 727
rect 2406 693 2436 710
rect 2406 676 2413 693
rect 2430 676 2436 693
rect 2406 659 2436 676
rect 2406 642 2413 659
rect 2430 642 2436 659
rect 2406 625 2436 642
rect 2406 608 2413 625
rect 2430 608 2436 625
rect 2406 591 2436 608
rect 2406 574 2413 591
rect 2430 574 2436 591
rect 2406 557 2436 574
rect 2406 540 2413 557
rect 2430 540 2436 557
rect 2406 523 2436 540
rect 2406 506 2413 523
rect 2430 506 2436 523
rect 2406 489 2436 506
rect 2406 472 2413 489
rect 2430 472 2436 489
rect 2406 455 2436 472
rect 2406 438 2413 455
rect 2430 438 2436 455
rect 2406 421 2436 438
rect 2406 404 2413 421
rect 2430 404 2436 421
rect 2406 387 2436 404
rect 2406 370 2413 387
rect 2430 370 2436 387
rect 2406 353 2436 370
rect 2406 336 2413 353
rect 2430 336 2436 353
rect 2406 319 2436 336
rect 2406 302 2413 319
rect 2430 302 2436 319
rect 2406 285 2436 302
rect 2406 268 2413 285
rect 2430 268 2436 285
rect 2406 251 2436 268
rect 2406 234 2413 251
rect 2430 234 2436 251
rect 2406 217 2436 234
rect 2406 200 2413 217
rect 2430 200 2436 217
rect 2406 183 2436 200
rect 2406 166 2413 183
rect 2430 166 2436 183
rect 2406 150 2436 166
rect 2451 1135 2482 1150
rect 2451 1118 2458 1135
rect 2475 1118 2482 1135
rect 2451 1101 2482 1118
rect 2451 1084 2458 1101
rect 2475 1084 2482 1101
rect 2451 1067 2482 1084
rect 2451 1050 2458 1067
rect 2475 1050 2482 1067
rect 2451 1033 2482 1050
rect 2451 1016 2458 1033
rect 2475 1016 2482 1033
rect 2451 999 2482 1016
rect 2451 982 2459 999
rect 2476 982 2482 999
rect 2451 965 2482 982
rect 2451 948 2459 965
rect 2476 948 2482 965
rect 2451 931 2482 948
rect 2451 914 2459 931
rect 2476 914 2482 931
rect 2451 897 2482 914
rect 2451 880 2459 897
rect 2476 880 2482 897
rect 2451 863 2482 880
rect 2451 846 2459 863
rect 2476 846 2482 863
rect 2451 829 2482 846
rect 2451 812 2459 829
rect 2476 812 2482 829
rect 2451 795 2482 812
rect 2451 778 2459 795
rect 2476 778 2482 795
rect 2451 761 2482 778
rect 2451 744 2459 761
rect 2476 744 2482 761
rect 2451 727 2482 744
rect 2451 710 2459 727
rect 2476 710 2482 727
rect 2451 693 2482 710
rect 2451 676 2459 693
rect 2476 676 2482 693
rect 2451 659 2482 676
rect 2451 642 2459 659
rect 2476 642 2482 659
rect 2451 625 2482 642
rect 2451 608 2459 625
rect 2476 608 2482 625
rect 2451 591 2482 608
rect 2451 574 2459 591
rect 2476 574 2482 591
rect 2451 557 2482 574
rect 2451 540 2459 557
rect 2476 540 2482 557
rect 2451 523 2482 540
rect 2451 506 2459 523
rect 2476 506 2482 523
rect 2451 489 2482 506
rect 2451 472 2459 489
rect 2476 472 2482 489
rect 2451 455 2482 472
rect 2451 438 2459 455
rect 2476 438 2482 455
rect 2451 421 2482 438
rect 2451 404 2459 421
rect 2476 404 2482 421
rect 2451 387 2482 404
rect 2451 370 2459 387
rect 2476 370 2482 387
rect 2451 353 2482 370
rect 2451 336 2459 353
rect 2476 336 2482 353
rect 2451 319 2482 336
rect 2451 302 2459 319
rect 2476 302 2482 319
rect 2451 285 2482 302
rect 2451 268 2459 285
rect 2476 268 2482 285
rect 2451 251 2482 268
rect 2451 234 2459 251
rect 2476 234 2482 251
rect 2451 217 2482 234
rect 2451 200 2459 217
rect 2476 200 2482 217
rect 2451 183 2482 200
rect 2451 166 2459 183
rect 2476 166 2482 183
rect 2451 150 2482 166
rect 2497 1137 2526 1150
rect 2497 1120 2503 1137
rect 2520 1120 2526 1137
rect 2497 1103 2526 1120
rect 2497 1086 2503 1103
rect 2520 1086 2526 1103
rect 2497 1069 2526 1086
rect 2497 1052 2503 1069
rect 2520 1052 2526 1069
rect 2497 1035 2526 1052
rect 2497 1018 2503 1035
rect 2520 1018 2526 1035
rect 2497 1001 2526 1018
rect 2497 984 2503 1001
rect 2520 984 2526 1001
rect 2497 967 2526 984
rect 2497 950 2503 967
rect 2520 950 2526 967
rect 2497 933 2526 950
rect 2497 916 2503 933
rect 2520 916 2526 933
rect 2497 899 2526 916
rect 2497 882 2503 899
rect 2520 882 2526 899
rect 2497 865 2526 882
rect 2497 848 2503 865
rect 2520 848 2526 865
rect 2497 831 2526 848
rect 2497 814 2503 831
rect 2520 814 2526 831
rect 2497 797 2526 814
rect 2497 780 2503 797
rect 2520 780 2526 797
rect 2497 763 2526 780
rect 2497 746 2503 763
rect 2520 746 2526 763
rect 2497 729 2526 746
rect 2497 712 2503 729
rect 2520 712 2526 729
rect 2497 695 2526 712
rect 2497 678 2503 695
rect 2520 678 2526 695
rect 2497 661 2526 678
rect 2497 644 2503 661
rect 2520 644 2526 661
rect 2497 627 2526 644
rect 2497 610 2503 627
rect 2520 610 2526 627
rect 2497 593 2526 610
rect 2497 576 2503 593
rect 2520 576 2526 593
rect 2497 559 2526 576
rect 2497 542 2503 559
rect 2520 542 2526 559
rect 2497 525 2526 542
rect 2497 508 2503 525
rect 2520 508 2526 525
rect 2497 491 2526 508
rect 2497 474 2503 491
rect 2520 474 2526 491
rect 2497 457 2526 474
rect 2497 440 2503 457
rect 2520 440 2526 457
rect 2497 423 2526 440
rect 2497 406 2503 423
rect 2520 406 2526 423
rect 2497 389 2526 406
rect 2497 372 2503 389
rect 2520 372 2526 389
rect 2497 355 2526 372
rect 2497 338 2503 355
rect 2520 338 2526 355
rect 2497 321 2526 338
rect 2497 304 2503 321
rect 2520 304 2526 321
rect 2497 287 2526 304
rect 2497 270 2503 287
rect 2520 270 2526 287
rect 2497 253 2526 270
rect 2497 236 2503 253
rect 2520 236 2526 253
rect 2497 219 2526 236
rect 2497 202 2503 219
rect 2520 202 2526 219
rect 2497 185 2526 202
rect 2497 168 2503 185
rect 2520 168 2526 185
rect 2497 150 2526 168
rect 2541 1135 2571 1150
rect 2541 1118 2547 1135
rect 2564 1118 2571 1135
rect 2541 1101 2571 1118
rect 2541 1084 2547 1101
rect 2564 1084 2571 1101
rect 2541 1067 2571 1084
rect 2541 1050 2547 1067
rect 2564 1050 2571 1067
rect 2541 1033 2571 1050
rect 2541 1016 2547 1033
rect 2564 1016 2571 1033
rect 2541 999 2571 1016
rect 2541 982 2548 999
rect 2565 982 2571 999
rect 2541 965 2571 982
rect 2541 948 2548 965
rect 2565 948 2571 965
rect 2541 931 2571 948
rect 2541 914 2548 931
rect 2565 914 2571 931
rect 2541 897 2571 914
rect 2541 880 2548 897
rect 2565 880 2571 897
rect 2541 863 2571 880
rect 2541 846 2548 863
rect 2565 846 2571 863
rect 2541 829 2571 846
rect 2541 812 2548 829
rect 2565 812 2571 829
rect 2541 795 2571 812
rect 2541 778 2548 795
rect 2565 778 2571 795
rect 2541 761 2571 778
rect 2541 744 2548 761
rect 2565 744 2571 761
rect 2541 727 2571 744
rect 2541 710 2548 727
rect 2565 710 2571 727
rect 2541 693 2571 710
rect 2541 676 2548 693
rect 2565 676 2571 693
rect 2541 659 2571 676
rect 2541 642 2548 659
rect 2565 642 2571 659
rect 2541 625 2571 642
rect 2541 608 2548 625
rect 2565 608 2571 625
rect 2541 591 2571 608
rect 2541 574 2548 591
rect 2565 574 2571 591
rect 2541 557 2571 574
rect 2541 540 2548 557
rect 2565 540 2571 557
rect 2541 523 2571 540
rect 2541 506 2548 523
rect 2565 506 2571 523
rect 2541 489 2571 506
rect 2541 472 2548 489
rect 2565 472 2571 489
rect 2541 455 2571 472
rect 2541 438 2548 455
rect 2565 438 2571 455
rect 2541 421 2571 438
rect 2541 404 2548 421
rect 2565 404 2571 421
rect 2541 387 2571 404
rect 2541 370 2548 387
rect 2565 370 2571 387
rect 2541 353 2571 370
rect 2541 336 2548 353
rect 2565 336 2571 353
rect 2541 319 2571 336
rect 2541 302 2548 319
rect 2565 302 2571 319
rect 2541 285 2571 302
rect 2541 268 2548 285
rect 2565 268 2571 285
rect 2541 251 2571 268
rect 2541 234 2548 251
rect 2565 234 2571 251
rect 2541 217 2571 234
rect 2541 200 2548 217
rect 2565 200 2571 217
rect 2541 183 2571 200
rect 2541 166 2548 183
rect 2565 166 2571 183
rect 2541 150 2571 166
rect 2586 1135 2616 1150
rect 2586 1118 2592 1135
rect 2609 1118 2616 1135
rect 2586 1101 2616 1118
rect 2586 1084 2592 1101
rect 2609 1084 2616 1101
rect 2586 1067 2616 1084
rect 2586 1050 2592 1067
rect 2609 1050 2616 1067
rect 2586 1033 2616 1050
rect 2586 1016 2592 1033
rect 2609 1016 2616 1033
rect 2586 999 2616 1016
rect 2586 982 2593 999
rect 2610 982 2616 999
rect 2586 965 2616 982
rect 2586 948 2593 965
rect 2610 948 2616 965
rect 2586 931 2616 948
rect 2586 914 2593 931
rect 2610 914 2616 931
rect 2586 897 2616 914
rect 2586 880 2593 897
rect 2610 880 2616 897
rect 2586 863 2616 880
rect 2586 846 2593 863
rect 2610 846 2616 863
rect 2586 829 2616 846
rect 2586 812 2593 829
rect 2610 812 2616 829
rect 2586 795 2616 812
rect 2586 778 2593 795
rect 2610 778 2616 795
rect 2586 761 2616 778
rect 2586 744 2593 761
rect 2610 744 2616 761
rect 2586 727 2616 744
rect 2586 710 2593 727
rect 2610 710 2616 727
rect 2586 693 2616 710
rect 2586 676 2593 693
rect 2610 676 2616 693
rect 2586 659 2616 676
rect 2586 642 2593 659
rect 2610 642 2616 659
rect 2586 625 2616 642
rect 2586 608 2593 625
rect 2610 608 2616 625
rect 2586 591 2616 608
rect 2586 574 2593 591
rect 2610 574 2616 591
rect 2586 557 2616 574
rect 2586 540 2593 557
rect 2610 540 2616 557
rect 2586 523 2616 540
rect 2586 506 2593 523
rect 2610 506 2616 523
rect 2586 489 2616 506
rect 2586 472 2593 489
rect 2610 472 2616 489
rect 2586 455 2616 472
rect 2586 438 2593 455
rect 2610 438 2616 455
rect 2586 421 2616 438
rect 2586 404 2593 421
rect 2610 404 2616 421
rect 2586 387 2616 404
rect 2586 370 2593 387
rect 2610 370 2616 387
rect 2586 353 2616 370
rect 2586 336 2593 353
rect 2610 336 2616 353
rect 2586 319 2616 336
rect 2586 302 2593 319
rect 2610 302 2616 319
rect 2586 285 2616 302
rect 2586 268 2593 285
rect 2610 268 2616 285
rect 2586 251 2616 268
rect 2586 234 2593 251
rect 2610 234 2616 251
rect 2586 217 2616 234
rect 2586 200 2593 217
rect 2610 200 2616 217
rect 2586 183 2616 200
rect 2586 166 2593 183
rect 2610 166 2616 183
rect 2586 150 2616 166
rect 2631 1135 2660 1150
rect 2631 1118 2637 1135
rect 2654 1118 2660 1135
rect 2631 1101 2660 1118
rect 2631 1084 2637 1101
rect 2654 1084 2660 1101
rect 2631 1067 2660 1084
rect 2631 1050 2637 1067
rect 2654 1050 2660 1067
rect 2631 1033 2660 1050
rect 2631 1016 2637 1033
rect 2654 1016 2660 1033
rect 2631 999 2660 1016
rect 2631 982 2638 999
rect 2655 982 2660 999
rect 2631 965 2660 982
rect 2631 948 2638 965
rect 2655 948 2660 965
rect 2631 931 2660 948
rect 2631 914 2638 931
rect 2655 914 2660 931
rect 2631 897 2660 914
rect 2631 880 2638 897
rect 2655 880 2660 897
rect 2631 863 2660 880
rect 2631 846 2638 863
rect 2655 846 2660 863
rect 2631 829 2660 846
rect 2631 812 2638 829
rect 2655 812 2660 829
rect 2631 795 2660 812
rect 2631 778 2638 795
rect 2655 778 2660 795
rect 2631 761 2660 778
rect 2631 744 2638 761
rect 2655 744 2660 761
rect 2631 727 2660 744
rect 2631 710 2638 727
rect 2655 710 2660 727
rect 2631 693 2660 710
rect 2631 676 2638 693
rect 2655 676 2660 693
rect 2631 659 2660 676
rect 2631 642 2638 659
rect 2655 642 2660 659
rect 2631 625 2660 642
rect 2631 608 2638 625
rect 2655 608 2660 625
rect 2631 591 2660 608
rect 2631 574 2638 591
rect 2655 574 2660 591
rect 2631 557 2660 574
rect 2631 540 2638 557
rect 2655 540 2660 557
rect 2631 523 2660 540
rect 2631 506 2638 523
rect 2655 506 2660 523
rect 2631 489 2660 506
rect 2631 472 2638 489
rect 2655 472 2660 489
rect 2631 455 2660 472
rect 2631 438 2638 455
rect 2655 438 2660 455
rect 2631 421 2660 438
rect 2631 404 2638 421
rect 2655 404 2660 421
rect 2631 387 2660 404
rect 2631 370 2638 387
rect 2655 370 2660 387
rect 2631 353 2660 370
rect 2631 336 2638 353
rect 2655 336 2660 353
rect 2631 319 2660 336
rect 2631 302 2638 319
rect 2655 302 2660 319
rect 2631 285 2660 302
rect 2631 268 2638 285
rect 2655 268 2660 285
rect 2631 251 2660 268
rect 2631 234 2638 251
rect 2655 234 2660 251
rect 2631 217 2660 234
rect 2631 200 2638 217
rect 2655 200 2660 217
rect 2631 183 2660 200
rect 2631 166 2638 183
rect 2655 166 2660 183
rect 2631 150 2660 166
<< ndiffc >>
rect -59 1118 -42 1135
rect -59 1084 -42 1101
rect -59 1050 -42 1067
rect -59 1016 -42 1033
rect -58 982 -41 999
rect -58 948 -41 965
rect -58 914 -41 931
rect -58 880 -41 897
rect -58 846 -41 863
rect -58 812 -41 829
rect -58 778 -41 795
rect -58 744 -41 761
rect -58 710 -41 727
rect -58 676 -41 693
rect -58 642 -41 659
rect -58 608 -41 625
rect -58 574 -41 591
rect -58 540 -41 557
rect -58 506 -41 523
rect -58 472 -41 489
rect -58 438 -41 455
rect -58 404 -41 421
rect -58 370 -41 387
rect -58 336 -41 353
rect -58 302 -41 319
rect -58 268 -41 285
rect -58 234 -41 251
rect -58 200 -41 217
rect -58 166 -41 183
rect -14 1120 3 1137
rect -14 1086 3 1103
rect -14 1052 3 1069
rect -14 1018 3 1035
rect -14 984 3 1001
rect -14 950 3 967
rect -14 916 3 933
rect -14 882 3 899
rect -14 848 3 865
rect -14 814 3 831
rect -14 780 3 797
rect -14 746 3 763
rect -14 712 3 729
rect -14 678 3 695
rect -14 644 3 661
rect -14 610 3 627
rect -14 576 3 593
rect -14 542 3 559
rect -14 508 3 525
rect -14 474 3 491
rect -14 440 3 457
rect -14 406 3 423
rect -14 372 3 389
rect -14 338 3 355
rect -14 304 3 321
rect -14 270 3 287
rect -14 236 3 253
rect -14 202 3 219
rect -14 168 3 185
rect 30 1118 47 1135
rect 30 1084 47 1101
rect 30 1050 47 1067
rect 30 1016 47 1033
rect 31 982 48 999
rect 31 948 48 965
rect 31 914 48 931
rect 31 880 48 897
rect 31 846 48 863
rect 31 812 48 829
rect 31 778 48 795
rect 31 744 48 761
rect 31 710 48 727
rect 31 676 48 693
rect 31 642 48 659
rect 31 608 48 625
rect 31 574 48 591
rect 31 540 48 557
rect 31 506 48 523
rect 31 472 48 489
rect 31 438 48 455
rect 31 404 48 421
rect 31 370 48 387
rect 31 336 48 353
rect 31 302 48 319
rect 31 268 48 285
rect 31 234 48 251
rect 31 200 48 217
rect 31 166 48 183
rect 75 1118 92 1135
rect 75 1084 92 1101
rect 75 1050 92 1067
rect 75 1016 92 1033
rect 76 982 93 999
rect 76 948 93 965
rect 76 914 93 931
rect 76 880 93 897
rect 76 846 93 863
rect 76 812 93 829
rect 76 778 93 795
rect 76 744 93 761
rect 76 710 93 727
rect 76 676 93 693
rect 76 642 93 659
rect 76 608 93 625
rect 76 574 93 591
rect 76 540 93 557
rect 76 506 93 523
rect 76 472 93 489
rect 76 438 93 455
rect 76 404 93 421
rect 76 370 93 387
rect 76 336 93 353
rect 76 302 93 319
rect 76 268 93 285
rect 76 234 93 251
rect 76 200 93 217
rect 76 166 93 183
rect 120 1118 137 1135
rect 120 1084 137 1101
rect 120 1050 137 1067
rect 120 1016 137 1033
rect 121 982 138 999
rect 121 948 138 965
rect 121 914 138 931
rect 121 880 138 897
rect 121 846 138 863
rect 121 812 138 829
rect 121 778 138 795
rect 121 744 138 761
rect 121 710 138 727
rect 121 676 138 693
rect 121 642 138 659
rect 121 608 138 625
rect 121 574 138 591
rect 121 540 138 557
rect 121 506 138 523
rect 121 472 138 489
rect 121 438 138 455
rect 121 404 138 421
rect 121 370 138 387
rect 121 336 138 353
rect 121 302 138 319
rect 121 268 138 285
rect 121 234 138 251
rect 121 200 138 217
rect 121 166 138 183
rect 165 1118 182 1135
rect 165 1084 182 1101
rect 165 1050 182 1067
rect 165 1016 182 1033
rect 166 982 183 999
rect 166 948 183 965
rect 166 914 183 931
rect 166 880 183 897
rect 166 846 183 863
rect 166 812 183 829
rect 166 778 183 795
rect 166 744 183 761
rect 166 710 183 727
rect 166 676 183 693
rect 166 642 183 659
rect 166 608 183 625
rect 166 574 183 591
rect 166 540 183 557
rect 166 506 183 523
rect 166 472 183 489
rect 166 438 183 455
rect 166 404 183 421
rect 166 370 183 387
rect 166 336 183 353
rect 166 302 183 319
rect 166 268 183 285
rect 166 234 183 251
rect 166 200 183 217
rect 166 166 183 183
rect 210 1118 227 1135
rect 210 1084 227 1101
rect 210 1050 227 1067
rect 210 1016 227 1033
rect 211 982 228 999
rect 211 948 228 965
rect 211 914 228 931
rect 211 880 228 897
rect 211 846 228 863
rect 211 812 228 829
rect 211 778 228 795
rect 211 744 228 761
rect 211 710 228 727
rect 211 676 228 693
rect 211 642 228 659
rect 211 608 228 625
rect 211 574 228 591
rect 211 540 228 557
rect 211 506 228 523
rect 211 472 228 489
rect 211 438 228 455
rect 211 404 228 421
rect 211 370 228 387
rect 211 336 228 353
rect 211 302 228 319
rect 211 268 228 285
rect 211 234 228 251
rect 211 200 228 217
rect 211 166 228 183
rect 255 1118 272 1135
rect 255 1084 272 1101
rect 255 1050 272 1067
rect 255 1016 272 1033
rect 256 982 273 999
rect 256 948 273 965
rect 256 914 273 931
rect 256 880 273 897
rect 256 846 273 863
rect 256 812 273 829
rect 256 778 273 795
rect 256 744 273 761
rect 256 710 273 727
rect 256 676 273 693
rect 256 642 273 659
rect 256 608 273 625
rect 256 574 273 591
rect 256 540 273 557
rect 256 506 273 523
rect 256 472 273 489
rect 256 438 273 455
rect 256 404 273 421
rect 256 370 273 387
rect 256 336 273 353
rect 256 302 273 319
rect 256 268 273 285
rect 256 234 273 251
rect 256 200 273 217
rect 256 166 273 183
rect 301 1118 318 1135
rect 301 1084 318 1101
rect 301 1050 318 1067
rect 301 1016 318 1033
rect 302 982 319 999
rect 302 948 319 965
rect 302 914 319 931
rect 302 880 319 897
rect 302 846 319 863
rect 302 812 319 829
rect 302 778 319 795
rect 302 744 319 761
rect 302 710 319 727
rect 302 676 319 693
rect 302 642 319 659
rect 302 608 319 625
rect 302 574 319 591
rect 302 540 319 557
rect 302 506 319 523
rect 302 472 319 489
rect 302 438 319 455
rect 302 404 319 421
rect 302 370 319 387
rect 302 336 319 353
rect 302 302 319 319
rect 302 268 319 285
rect 302 234 319 251
rect 302 200 319 217
rect 302 166 319 183
rect 346 1120 363 1137
rect 346 1086 363 1103
rect 346 1052 363 1069
rect 346 1018 363 1035
rect 346 984 363 1001
rect 346 950 363 967
rect 346 916 363 933
rect 346 882 363 899
rect 346 848 363 865
rect 346 814 363 831
rect 346 780 363 797
rect 346 746 363 763
rect 346 712 363 729
rect 346 678 363 695
rect 346 644 363 661
rect 346 610 363 627
rect 346 576 363 593
rect 346 542 363 559
rect 346 508 363 525
rect 346 474 363 491
rect 346 440 363 457
rect 346 406 363 423
rect 346 372 363 389
rect 346 338 363 355
rect 346 304 363 321
rect 346 270 363 287
rect 346 236 363 253
rect 346 202 363 219
rect 346 168 363 185
rect 390 1118 407 1135
rect 390 1084 407 1101
rect 390 1050 407 1067
rect 390 1016 407 1033
rect 391 982 408 999
rect 391 948 408 965
rect 391 914 408 931
rect 391 880 408 897
rect 391 846 408 863
rect 391 812 408 829
rect 391 778 408 795
rect 391 744 408 761
rect 391 710 408 727
rect 391 676 408 693
rect 391 642 408 659
rect 391 608 408 625
rect 391 574 408 591
rect 391 540 408 557
rect 391 506 408 523
rect 391 472 408 489
rect 391 438 408 455
rect 391 404 408 421
rect 391 370 408 387
rect 391 336 408 353
rect 391 302 408 319
rect 391 268 408 285
rect 391 234 408 251
rect 391 200 408 217
rect 391 166 408 183
rect 435 1118 452 1135
rect 435 1084 452 1101
rect 435 1050 452 1067
rect 435 1016 452 1033
rect 436 982 453 999
rect 436 948 453 965
rect 436 914 453 931
rect 436 880 453 897
rect 436 846 453 863
rect 436 812 453 829
rect 436 778 453 795
rect 436 744 453 761
rect 436 710 453 727
rect 436 676 453 693
rect 436 642 453 659
rect 436 608 453 625
rect 436 574 453 591
rect 436 540 453 557
rect 436 506 453 523
rect 436 472 453 489
rect 436 438 453 455
rect 436 404 453 421
rect 436 370 453 387
rect 436 336 453 353
rect 436 302 453 319
rect 436 268 453 285
rect 436 234 453 251
rect 436 200 453 217
rect 436 166 453 183
rect 480 1118 497 1135
rect 480 1084 497 1101
rect 480 1050 497 1067
rect 480 1016 497 1033
rect 481 982 498 999
rect 481 948 498 965
rect 481 914 498 931
rect 481 880 498 897
rect 481 846 498 863
rect 481 812 498 829
rect 481 778 498 795
rect 481 744 498 761
rect 481 710 498 727
rect 481 676 498 693
rect 481 642 498 659
rect 481 608 498 625
rect 481 574 498 591
rect 481 540 498 557
rect 481 506 498 523
rect 481 472 498 489
rect 481 438 498 455
rect 481 404 498 421
rect 481 370 498 387
rect 481 336 498 353
rect 481 302 498 319
rect 481 268 498 285
rect 481 234 498 251
rect 481 200 498 217
rect 481 166 498 183
rect 525 1118 542 1135
rect 525 1084 542 1101
rect 525 1050 542 1067
rect 525 1016 542 1033
rect 526 982 543 999
rect 526 948 543 965
rect 526 914 543 931
rect 526 880 543 897
rect 526 846 543 863
rect 526 812 543 829
rect 526 778 543 795
rect 526 744 543 761
rect 526 710 543 727
rect 526 676 543 693
rect 526 642 543 659
rect 526 608 543 625
rect 526 574 543 591
rect 526 540 543 557
rect 526 506 543 523
rect 526 472 543 489
rect 526 438 543 455
rect 526 404 543 421
rect 526 370 543 387
rect 526 336 543 353
rect 526 302 543 319
rect 526 268 543 285
rect 526 234 543 251
rect 526 200 543 217
rect 526 166 543 183
rect 570 1118 587 1135
rect 570 1084 587 1101
rect 570 1050 587 1067
rect 570 1016 587 1033
rect 571 982 588 999
rect 571 948 588 965
rect 571 914 588 931
rect 571 880 588 897
rect 571 846 588 863
rect 571 812 588 829
rect 571 778 588 795
rect 571 744 588 761
rect 571 710 588 727
rect 571 676 588 693
rect 571 642 588 659
rect 571 608 588 625
rect 571 574 588 591
rect 571 540 588 557
rect 571 506 588 523
rect 571 472 588 489
rect 571 438 588 455
rect 571 404 588 421
rect 571 370 588 387
rect 571 336 588 353
rect 571 302 588 319
rect 571 268 588 285
rect 571 234 588 251
rect 571 200 588 217
rect 571 166 588 183
rect 615 1118 632 1135
rect 615 1084 632 1101
rect 615 1050 632 1067
rect 615 1016 632 1033
rect 616 982 633 999
rect 616 948 633 965
rect 616 914 633 931
rect 616 880 633 897
rect 616 846 633 863
rect 616 812 633 829
rect 616 778 633 795
rect 616 744 633 761
rect 616 710 633 727
rect 616 676 633 693
rect 616 642 633 659
rect 616 608 633 625
rect 616 574 633 591
rect 616 540 633 557
rect 616 506 633 523
rect 616 472 633 489
rect 616 438 633 455
rect 616 404 633 421
rect 616 370 633 387
rect 616 336 633 353
rect 616 302 633 319
rect 616 268 633 285
rect 616 234 633 251
rect 616 200 633 217
rect 616 166 633 183
rect 660 1118 677 1135
rect 660 1084 677 1101
rect 660 1050 677 1067
rect 660 1016 677 1033
rect 661 982 678 999
rect 661 948 678 965
rect 661 914 678 931
rect 661 880 678 897
rect 661 846 678 863
rect 661 812 678 829
rect 661 778 678 795
rect 661 744 678 761
rect 661 710 678 727
rect 661 676 678 693
rect 661 642 678 659
rect 661 608 678 625
rect 661 574 678 591
rect 661 540 678 557
rect 661 506 678 523
rect 661 472 678 489
rect 661 438 678 455
rect 661 404 678 421
rect 661 370 678 387
rect 661 336 678 353
rect 661 302 678 319
rect 661 268 678 285
rect 661 234 678 251
rect 661 200 678 217
rect 661 166 678 183
rect 705 1120 722 1137
rect 705 1086 722 1103
rect 705 1052 722 1069
rect 705 1018 722 1035
rect 705 984 722 1001
rect 705 950 722 967
rect 705 916 722 933
rect 705 882 722 899
rect 705 848 722 865
rect 705 814 722 831
rect 705 780 722 797
rect 705 746 722 763
rect 705 712 722 729
rect 705 678 722 695
rect 705 644 722 661
rect 705 610 722 627
rect 705 576 722 593
rect 705 542 722 559
rect 705 508 722 525
rect 705 474 722 491
rect 705 440 722 457
rect 705 406 722 423
rect 705 372 722 389
rect 705 338 722 355
rect 705 304 722 321
rect 705 270 722 287
rect 705 236 722 253
rect 705 202 722 219
rect 705 168 722 185
rect 749 1118 766 1135
rect 749 1084 766 1101
rect 749 1050 766 1067
rect 749 1016 766 1033
rect 750 982 767 999
rect 750 948 767 965
rect 750 914 767 931
rect 750 880 767 897
rect 750 846 767 863
rect 750 812 767 829
rect 750 778 767 795
rect 750 744 767 761
rect 750 710 767 727
rect 750 676 767 693
rect 750 642 767 659
rect 750 608 767 625
rect 750 574 767 591
rect 750 540 767 557
rect 750 506 767 523
rect 750 472 767 489
rect 750 438 767 455
rect 750 404 767 421
rect 750 370 767 387
rect 750 336 767 353
rect 750 302 767 319
rect 750 268 767 285
rect 750 234 767 251
rect 750 200 767 217
rect 750 166 767 183
rect 794 1118 811 1135
rect 794 1084 811 1101
rect 794 1050 811 1067
rect 794 1016 811 1033
rect 795 982 812 999
rect 795 948 812 965
rect 795 914 812 931
rect 795 880 812 897
rect 795 846 812 863
rect 795 812 812 829
rect 795 778 812 795
rect 795 744 812 761
rect 795 710 812 727
rect 795 676 812 693
rect 795 642 812 659
rect 795 608 812 625
rect 795 574 812 591
rect 795 540 812 557
rect 795 506 812 523
rect 795 472 812 489
rect 795 438 812 455
rect 795 404 812 421
rect 795 370 812 387
rect 795 336 812 353
rect 795 302 812 319
rect 795 268 812 285
rect 795 234 812 251
rect 795 200 812 217
rect 795 166 812 183
rect 839 1118 856 1135
rect 839 1084 856 1101
rect 839 1050 856 1067
rect 839 1016 856 1033
rect 840 982 857 999
rect 840 948 857 965
rect 840 914 857 931
rect 840 880 857 897
rect 840 846 857 863
rect 840 812 857 829
rect 840 778 857 795
rect 840 744 857 761
rect 840 710 857 727
rect 840 676 857 693
rect 840 642 857 659
rect 840 608 857 625
rect 840 574 857 591
rect 840 540 857 557
rect 840 506 857 523
rect 840 472 857 489
rect 840 438 857 455
rect 840 404 857 421
rect 840 370 857 387
rect 840 336 857 353
rect 840 302 857 319
rect 840 268 857 285
rect 840 234 857 251
rect 840 200 857 217
rect 840 166 857 183
rect 884 1118 901 1135
rect 884 1084 901 1101
rect 884 1050 901 1067
rect 884 1016 901 1033
rect 885 982 902 999
rect 885 948 902 965
rect 885 914 902 931
rect 885 880 902 897
rect 885 846 902 863
rect 885 812 902 829
rect 885 778 902 795
rect 885 744 902 761
rect 885 710 902 727
rect 885 676 902 693
rect 885 642 902 659
rect 885 608 902 625
rect 885 574 902 591
rect 885 540 902 557
rect 885 506 902 523
rect 885 472 902 489
rect 885 438 902 455
rect 885 404 902 421
rect 885 370 902 387
rect 885 336 902 353
rect 885 302 902 319
rect 885 268 902 285
rect 885 234 902 251
rect 885 200 902 217
rect 885 166 902 183
rect 929 1118 946 1135
rect 929 1084 946 1101
rect 929 1050 946 1067
rect 929 1016 946 1033
rect 930 982 947 999
rect 930 948 947 965
rect 930 914 947 931
rect 930 880 947 897
rect 930 846 947 863
rect 930 812 947 829
rect 930 778 947 795
rect 930 744 947 761
rect 930 710 947 727
rect 930 676 947 693
rect 930 642 947 659
rect 930 608 947 625
rect 930 574 947 591
rect 930 540 947 557
rect 930 506 947 523
rect 930 472 947 489
rect 930 438 947 455
rect 930 404 947 421
rect 930 370 947 387
rect 930 336 947 353
rect 930 302 947 319
rect 930 268 947 285
rect 930 234 947 251
rect 930 200 947 217
rect 930 166 947 183
rect 974 1118 991 1135
rect 974 1084 991 1101
rect 974 1050 991 1067
rect 974 1016 991 1033
rect 975 982 992 999
rect 975 948 992 965
rect 975 914 992 931
rect 975 880 992 897
rect 975 846 992 863
rect 975 812 992 829
rect 975 778 992 795
rect 975 744 992 761
rect 975 710 992 727
rect 975 676 992 693
rect 975 642 992 659
rect 975 608 992 625
rect 975 574 992 591
rect 975 540 992 557
rect 975 506 992 523
rect 975 472 992 489
rect 975 438 992 455
rect 975 404 992 421
rect 975 370 992 387
rect 975 336 992 353
rect 975 302 992 319
rect 975 268 992 285
rect 975 234 992 251
rect 975 200 992 217
rect 975 166 992 183
rect 1020 1118 1037 1135
rect 1020 1084 1037 1101
rect 1020 1050 1037 1067
rect 1020 1016 1037 1033
rect 1021 982 1038 999
rect 1021 948 1038 965
rect 1021 914 1038 931
rect 1021 880 1038 897
rect 1021 846 1038 863
rect 1021 812 1038 829
rect 1021 778 1038 795
rect 1021 744 1038 761
rect 1021 710 1038 727
rect 1021 676 1038 693
rect 1021 642 1038 659
rect 1021 608 1038 625
rect 1021 574 1038 591
rect 1021 540 1038 557
rect 1021 506 1038 523
rect 1021 472 1038 489
rect 1021 438 1038 455
rect 1021 404 1038 421
rect 1021 370 1038 387
rect 1021 336 1038 353
rect 1021 302 1038 319
rect 1021 268 1038 285
rect 1021 234 1038 251
rect 1021 200 1038 217
rect 1021 166 1038 183
rect 1065 1120 1082 1137
rect 1065 1086 1082 1103
rect 1065 1052 1082 1069
rect 1065 1018 1082 1035
rect 1065 984 1082 1001
rect 1065 950 1082 967
rect 1065 916 1082 933
rect 1065 882 1082 899
rect 1065 848 1082 865
rect 1065 814 1082 831
rect 1065 780 1082 797
rect 1065 746 1082 763
rect 1065 712 1082 729
rect 1065 678 1082 695
rect 1065 644 1082 661
rect 1065 610 1082 627
rect 1065 576 1082 593
rect 1065 542 1082 559
rect 1065 508 1082 525
rect 1065 474 1082 491
rect 1065 440 1082 457
rect 1065 406 1082 423
rect 1065 372 1082 389
rect 1065 338 1082 355
rect 1065 304 1082 321
rect 1065 270 1082 287
rect 1065 236 1082 253
rect 1065 202 1082 219
rect 1065 168 1082 185
rect 1109 1118 1126 1135
rect 1109 1084 1126 1101
rect 1109 1050 1126 1067
rect 1109 1016 1126 1033
rect 1110 982 1127 999
rect 1110 948 1127 965
rect 1110 914 1127 931
rect 1110 880 1127 897
rect 1110 846 1127 863
rect 1110 812 1127 829
rect 1110 778 1127 795
rect 1110 744 1127 761
rect 1110 710 1127 727
rect 1110 676 1127 693
rect 1110 642 1127 659
rect 1110 608 1127 625
rect 1110 574 1127 591
rect 1110 540 1127 557
rect 1110 506 1127 523
rect 1110 472 1127 489
rect 1110 438 1127 455
rect 1110 404 1127 421
rect 1110 370 1127 387
rect 1110 336 1127 353
rect 1110 302 1127 319
rect 1110 268 1127 285
rect 1110 234 1127 251
rect 1110 200 1127 217
rect 1110 166 1127 183
rect 1154 1118 1171 1135
rect 1154 1084 1171 1101
rect 1154 1050 1171 1067
rect 1154 1016 1171 1033
rect 1155 982 1172 999
rect 1155 948 1172 965
rect 1155 914 1172 931
rect 1155 880 1172 897
rect 1155 846 1172 863
rect 1155 812 1172 829
rect 1155 778 1172 795
rect 1155 744 1172 761
rect 1155 710 1172 727
rect 1155 676 1172 693
rect 1155 642 1172 659
rect 1155 608 1172 625
rect 1155 574 1172 591
rect 1155 540 1172 557
rect 1155 506 1172 523
rect 1155 472 1172 489
rect 1155 438 1172 455
rect 1155 404 1172 421
rect 1155 370 1172 387
rect 1155 336 1172 353
rect 1155 302 1172 319
rect 1155 268 1172 285
rect 1155 234 1172 251
rect 1155 200 1172 217
rect 1155 166 1172 183
rect 1199 1118 1216 1135
rect 1199 1084 1216 1101
rect 1199 1050 1216 1067
rect 1199 1016 1216 1033
rect 1200 982 1217 999
rect 1200 948 1217 965
rect 1200 914 1217 931
rect 1200 880 1217 897
rect 1200 846 1217 863
rect 1200 812 1217 829
rect 1200 778 1217 795
rect 1200 744 1217 761
rect 1200 710 1217 727
rect 1200 676 1217 693
rect 1200 642 1217 659
rect 1200 608 1217 625
rect 1200 574 1217 591
rect 1200 540 1217 557
rect 1200 506 1217 523
rect 1200 472 1217 489
rect 1200 438 1217 455
rect 1200 404 1217 421
rect 1200 370 1217 387
rect 1200 336 1217 353
rect 1200 302 1217 319
rect 1200 268 1217 285
rect 1200 234 1217 251
rect 1200 200 1217 217
rect 1200 166 1217 183
rect 1244 1118 1261 1135
rect 1244 1084 1261 1101
rect 1244 1050 1261 1067
rect 1244 1016 1261 1033
rect 1245 982 1262 999
rect 1245 948 1262 965
rect 1245 914 1262 931
rect 1245 880 1262 897
rect 1245 846 1262 863
rect 1245 812 1262 829
rect 1245 778 1262 795
rect 1245 744 1262 761
rect 1245 710 1262 727
rect 1245 676 1262 693
rect 1245 642 1262 659
rect 1245 608 1262 625
rect 1245 574 1262 591
rect 1245 540 1262 557
rect 1245 506 1262 523
rect 1245 472 1262 489
rect 1245 438 1262 455
rect 1245 404 1262 421
rect 1245 370 1262 387
rect 1245 336 1262 353
rect 1245 302 1262 319
rect 1245 268 1262 285
rect 1245 234 1262 251
rect 1245 200 1262 217
rect 1245 166 1262 183
rect 1289 1118 1306 1135
rect 1289 1084 1306 1101
rect 1289 1050 1306 1067
rect 1289 1016 1306 1033
rect 1290 982 1307 999
rect 1290 948 1307 965
rect 1290 914 1307 931
rect 1290 880 1307 897
rect 1290 846 1307 863
rect 1290 812 1307 829
rect 1290 778 1307 795
rect 1290 744 1307 761
rect 1290 710 1307 727
rect 1290 676 1307 693
rect 1290 642 1307 659
rect 1290 608 1307 625
rect 1290 574 1307 591
rect 1290 540 1307 557
rect 1290 506 1307 523
rect 1290 472 1307 489
rect 1290 438 1307 455
rect 1290 404 1307 421
rect 1290 370 1307 387
rect 1290 336 1307 353
rect 1290 302 1307 319
rect 1290 268 1307 285
rect 1290 234 1307 251
rect 1290 200 1307 217
rect 1290 166 1307 183
rect 1334 1118 1351 1135
rect 1334 1084 1351 1101
rect 1334 1050 1351 1067
rect 1334 1016 1351 1033
rect 1335 982 1352 999
rect 1335 948 1352 965
rect 1335 914 1352 931
rect 1335 880 1352 897
rect 1335 846 1352 863
rect 1335 812 1352 829
rect 1335 778 1352 795
rect 1335 744 1352 761
rect 1335 710 1352 727
rect 1335 676 1352 693
rect 1335 642 1352 659
rect 1335 608 1352 625
rect 1335 574 1352 591
rect 1335 540 1352 557
rect 1335 506 1352 523
rect 1335 472 1352 489
rect 1335 438 1352 455
rect 1335 404 1352 421
rect 1335 370 1352 387
rect 1335 336 1352 353
rect 1335 302 1352 319
rect 1335 268 1352 285
rect 1335 234 1352 251
rect 1335 200 1352 217
rect 1335 166 1352 183
rect 1379 1118 1396 1135
rect 1379 1084 1396 1101
rect 1379 1050 1396 1067
rect 1379 1016 1396 1033
rect 1380 982 1397 999
rect 1380 948 1397 965
rect 1380 914 1397 931
rect 1380 880 1397 897
rect 1380 846 1397 863
rect 1380 812 1397 829
rect 1380 778 1397 795
rect 1380 744 1397 761
rect 1380 710 1397 727
rect 1380 676 1397 693
rect 1380 642 1397 659
rect 1380 608 1397 625
rect 1380 574 1397 591
rect 1380 540 1397 557
rect 1380 506 1397 523
rect 1380 472 1397 489
rect 1380 438 1397 455
rect 1380 404 1397 421
rect 1380 370 1397 387
rect 1380 336 1397 353
rect 1380 302 1397 319
rect 1380 268 1397 285
rect 1380 234 1397 251
rect 1380 200 1397 217
rect 1380 166 1397 183
rect 1424 1120 1441 1137
rect 1424 1086 1441 1103
rect 1424 1052 1441 1069
rect 1424 1018 1441 1035
rect 1424 984 1441 1001
rect 1424 950 1441 967
rect 1424 916 1441 933
rect 1424 882 1441 899
rect 1424 848 1441 865
rect 1424 814 1441 831
rect 1424 780 1441 797
rect 1424 746 1441 763
rect 1424 712 1441 729
rect 1424 678 1441 695
rect 1424 644 1441 661
rect 1424 610 1441 627
rect 1424 576 1441 593
rect 1424 542 1441 559
rect 1424 508 1441 525
rect 1424 474 1441 491
rect 1424 440 1441 457
rect 1424 406 1441 423
rect 1424 372 1441 389
rect 1424 338 1441 355
rect 1424 304 1441 321
rect 1424 270 1441 287
rect 1424 236 1441 253
rect 1424 202 1441 219
rect 1424 168 1441 185
rect 1468 1118 1485 1135
rect 1468 1084 1485 1101
rect 1468 1050 1485 1067
rect 1468 1016 1485 1033
rect 1469 982 1486 999
rect 1469 948 1486 965
rect 1469 914 1486 931
rect 1469 880 1486 897
rect 1469 846 1486 863
rect 1469 812 1486 829
rect 1469 778 1486 795
rect 1469 744 1486 761
rect 1469 710 1486 727
rect 1469 676 1486 693
rect 1469 642 1486 659
rect 1469 608 1486 625
rect 1469 574 1486 591
rect 1469 540 1486 557
rect 1469 506 1486 523
rect 1469 472 1486 489
rect 1469 438 1486 455
rect 1469 404 1486 421
rect 1469 370 1486 387
rect 1469 336 1486 353
rect 1469 302 1486 319
rect 1469 268 1486 285
rect 1469 234 1486 251
rect 1469 200 1486 217
rect 1469 166 1486 183
rect 1513 1118 1530 1135
rect 1513 1084 1530 1101
rect 1513 1050 1530 1067
rect 1513 1016 1530 1033
rect 1514 982 1531 999
rect 1514 948 1531 965
rect 1514 914 1531 931
rect 1514 880 1531 897
rect 1514 846 1531 863
rect 1514 812 1531 829
rect 1514 778 1531 795
rect 1514 744 1531 761
rect 1514 710 1531 727
rect 1514 676 1531 693
rect 1514 642 1531 659
rect 1514 608 1531 625
rect 1514 574 1531 591
rect 1514 540 1531 557
rect 1514 506 1531 523
rect 1514 472 1531 489
rect 1514 438 1531 455
rect 1514 404 1531 421
rect 1514 370 1531 387
rect 1514 336 1531 353
rect 1514 302 1531 319
rect 1514 268 1531 285
rect 1514 234 1531 251
rect 1514 200 1531 217
rect 1514 166 1531 183
rect 1558 1118 1575 1135
rect 1558 1084 1575 1101
rect 1558 1050 1575 1067
rect 1558 1016 1575 1033
rect 1559 982 1576 999
rect 1559 948 1576 965
rect 1559 914 1576 931
rect 1559 880 1576 897
rect 1559 846 1576 863
rect 1559 812 1576 829
rect 1559 778 1576 795
rect 1559 744 1576 761
rect 1559 710 1576 727
rect 1559 676 1576 693
rect 1559 642 1576 659
rect 1559 608 1576 625
rect 1559 574 1576 591
rect 1559 540 1576 557
rect 1559 506 1576 523
rect 1559 472 1576 489
rect 1559 438 1576 455
rect 1559 404 1576 421
rect 1559 370 1576 387
rect 1559 336 1576 353
rect 1559 302 1576 319
rect 1559 268 1576 285
rect 1559 234 1576 251
rect 1559 200 1576 217
rect 1559 166 1576 183
rect 1603 1118 1620 1135
rect 1603 1084 1620 1101
rect 1603 1050 1620 1067
rect 1603 1016 1620 1033
rect 1604 982 1621 999
rect 1604 948 1621 965
rect 1604 914 1621 931
rect 1604 880 1621 897
rect 1604 846 1621 863
rect 1604 812 1621 829
rect 1604 778 1621 795
rect 1604 744 1621 761
rect 1604 710 1621 727
rect 1604 676 1621 693
rect 1604 642 1621 659
rect 1604 608 1621 625
rect 1604 574 1621 591
rect 1604 540 1621 557
rect 1604 506 1621 523
rect 1604 472 1621 489
rect 1604 438 1621 455
rect 1604 404 1621 421
rect 1604 370 1621 387
rect 1604 336 1621 353
rect 1604 302 1621 319
rect 1604 268 1621 285
rect 1604 234 1621 251
rect 1604 200 1621 217
rect 1604 166 1621 183
rect 1648 1118 1665 1135
rect 1648 1084 1665 1101
rect 1648 1050 1665 1067
rect 1648 1016 1665 1033
rect 1649 982 1666 999
rect 1649 948 1666 965
rect 1649 914 1666 931
rect 1649 880 1666 897
rect 1649 846 1666 863
rect 1649 812 1666 829
rect 1649 778 1666 795
rect 1649 744 1666 761
rect 1649 710 1666 727
rect 1649 676 1666 693
rect 1649 642 1666 659
rect 1649 608 1666 625
rect 1649 574 1666 591
rect 1649 540 1666 557
rect 1649 506 1666 523
rect 1649 472 1666 489
rect 1649 438 1666 455
rect 1649 404 1666 421
rect 1649 370 1666 387
rect 1649 336 1666 353
rect 1649 302 1666 319
rect 1649 268 1666 285
rect 1649 234 1666 251
rect 1649 200 1666 217
rect 1649 166 1666 183
rect 1693 1118 1710 1135
rect 1693 1084 1710 1101
rect 1693 1050 1710 1067
rect 1693 1016 1710 1033
rect 1694 982 1711 999
rect 1694 948 1711 965
rect 1694 914 1711 931
rect 1694 880 1711 897
rect 1694 846 1711 863
rect 1694 812 1711 829
rect 1694 778 1711 795
rect 1694 744 1711 761
rect 1694 710 1711 727
rect 1694 676 1711 693
rect 1694 642 1711 659
rect 1694 608 1711 625
rect 1694 574 1711 591
rect 1694 540 1711 557
rect 1694 506 1711 523
rect 1694 472 1711 489
rect 1694 438 1711 455
rect 1694 404 1711 421
rect 1694 370 1711 387
rect 1694 336 1711 353
rect 1694 302 1711 319
rect 1694 268 1711 285
rect 1694 234 1711 251
rect 1694 200 1711 217
rect 1694 166 1711 183
rect 1739 1118 1756 1135
rect 1739 1084 1756 1101
rect 1739 1050 1756 1067
rect 1739 1016 1756 1033
rect 1740 982 1757 999
rect 1740 948 1757 965
rect 1740 914 1757 931
rect 1740 880 1757 897
rect 1740 846 1757 863
rect 1740 812 1757 829
rect 1740 778 1757 795
rect 1740 744 1757 761
rect 1740 710 1757 727
rect 1740 676 1757 693
rect 1740 642 1757 659
rect 1740 608 1757 625
rect 1740 574 1757 591
rect 1740 540 1757 557
rect 1740 506 1757 523
rect 1740 472 1757 489
rect 1740 438 1757 455
rect 1740 404 1757 421
rect 1740 370 1757 387
rect 1740 336 1757 353
rect 1740 302 1757 319
rect 1740 268 1757 285
rect 1740 234 1757 251
rect 1740 200 1757 217
rect 1740 166 1757 183
rect 1784 1120 1801 1137
rect 1784 1086 1801 1103
rect 1784 1052 1801 1069
rect 1784 1018 1801 1035
rect 1784 984 1801 1001
rect 1784 950 1801 967
rect 1784 916 1801 933
rect 1784 882 1801 899
rect 1784 848 1801 865
rect 1784 814 1801 831
rect 1784 780 1801 797
rect 1784 746 1801 763
rect 1784 712 1801 729
rect 1784 678 1801 695
rect 1784 644 1801 661
rect 1784 610 1801 627
rect 1784 576 1801 593
rect 1784 542 1801 559
rect 1784 508 1801 525
rect 1784 474 1801 491
rect 1784 440 1801 457
rect 1784 406 1801 423
rect 1784 372 1801 389
rect 1784 338 1801 355
rect 1784 304 1801 321
rect 1784 270 1801 287
rect 1784 236 1801 253
rect 1784 202 1801 219
rect 1784 168 1801 185
rect 1828 1118 1845 1135
rect 1828 1084 1845 1101
rect 1828 1050 1845 1067
rect 1828 1016 1845 1033
rect 1829 982 1846 999
rect 1829 948 1846 965
rect 1829 914 1846 931
rect 1829 880 1846 897
rect 1829 846 1846 863
rect 1829 812 1846 829
rect 1829 778 1846 795
rect 1829 744 1846 761
rect 1829 710 1846 727
rect 1829 676 1846 693
rect 1829 642 1846 659
rect 1829 608 1846 625
rect 1829 574 1846 591
rect 1829 540 1846 557
rect 1829 506 1846 523
rect 1829 472 1846 489
rect 1829 438 1846 455
rect 1829 404 1846 421
rect 1829 370 1846 387
rect 1829 336 1846 353
rect 1829 302 1846 319
rect 1829 268 1846 285
rect 1829 234 1846 251
rect 1829 200 1846 217
rect 1829 166 1846 183
rect 1873 1118 1890 1135
rect 1873 1084 1890 1101
rect 1873 1050 1890 1067
rect 1873 1016 1890 1033
rect 1874 982 1891 999
rect 1874 948 1891 965
rect 1874 914 1891 931
rect 1874 880 1891 897
rect 1874 846 1891 863
rect 1874 812 1891 829
rect 1874 778 1891 795
rect 1874 744 1891 761
rect 1874 710 1891 727
rect 1874 676 1891 693
rect 1874 642 1891 659
rect 1874 608 1891 625
rect 1874 574 1891 591
rect 1874 540 1891 557
rect 1874 506 1891 523
rect 1874 472 1891 489
rect 1874 438 1891 455
rect 1874 404 1891 421
rect 1874 370 1891 387
rect 1874 336 1891 353
rect 1874 302 1891 319
rect 1874 268 1891 285
rect 1874 234 1891 251
rect 1874 200 1891 217
rect 1874 166 1891 183
rect 1918 1118 1935 1135
rect 1918 1084 1935 1101
rect 1918 1050 1935 1067
rect 1918 1016 1935 1033
rect 1919 982 1936 999
rect 1919 948 1936 965
rect 1919 914 1936 931
rect 1919 880 1936 897
rect 1919 846 1936 863
rect 1919 812 1936 829
rect 1919 778 1936 795
rect 1919 744 1936 761
rect 1919 710 1936 727
rect 1919 676 1936 693
rect 1919 642 1936 659
rect 1919 608 1936 625
rect 1919 574 1936 591
rect 1919 540 1936 557
rect 1919 506 1936 523
rect 1919 472 1936 489
rect 1919 438 1936 455
rect 1919 404 1936 421
rect 1919 370 1936 387
rect 1919 336 1936 353
rect 1919 302 1936 319
rect 1919 268 1936 285
rect 1919 234 1936 251
rect 1919 200 1936 217
rect 1919 166 1936 183
rect 1963 1118 1980 1135
rect 1963 1084 1980 1101
rect 1963 1050 1980 1067
rect 1963 1016 1980 1033
rect 1964 982 1981 999
rect 1964 948 1981 965
rect 1964 914 1981 931
rect 1964 880 1981 897
rect 1964 846 1981 863
rect 1964 812 1981 829
rect 1964 778 1981 795
rect 1964 744 1981 761
rect 1964 710 1981 727
rect 1964 676 1981 693
rect 1964 642 1981 659
rect 1964 608 1981 625
rect 1964 574 1981 591
rect 1964 540 1981 557
rect 1964 506 1981 523
rect 1964 472 1981 489
rect 1964 438 1981 455
rect 1964 404 1981 421
rect 1964 370 1981 387
rect 1964 336 1981 353
rect 1964 302 1981 319
rect 1964 268 1981 285
rect 1964 234 1981 251
rect 1964 200 1981 217
rect 1964 166 1981 183
rect 2008 1118 2025 1135
rect 2008 1084 2025 1101
rect 2008 1050 2025 1067
rect 2008 1016 2025 1033
rect 2009 982 2026 999
rect 2009 948 2026 965
rect 2009 914 2026 931
rect 2009 880 2026 897
rect 2009 846 2026 863
rect 2009 812 2026 829
rect 2009 778 2026 795
rect 2009 744 2026 761
rect 2009 710 2026 727
rect 2009 676 2026 693
rect 2009 642 2026 659
rect 2009 608 2026 625
rect 2009 574 2026 591
rect 2009 540 2026 557
rect 2009 506 2026 523
rect 2009 472 2026 489
rect 2009 438 2026 455
rect 2009 404 2026 421
rect 2009 370 2026 387
rect 2009 336 2026 353
rect 2009 302 2026 319
rect 2009 268 2026 285
rect 2009 234 2026 251
rect 2009 200 2026 217
rect 2009 166 2026 183
rect 2053 1118 2070 1135
rect 2053 1084 2070 1101
rect 2053 1050 2070 1067
rect 2053 1016 2070 1033
rect 2054 982 2071 999
rect 2054 948 2071 965
rect 2054 914 2071 931
rect 2054 880 2071 897
rect 2054 846 2071 863
rect 2054 812 2071 829
rect 2054 778 2071 795
rect 2054 744 2071 761
rect 2054 710 2071 727
rect 2054 676 2071 693
rect 2054 642 2071 659
rect 2054 608 2071 625
rect 2054 574 2071 591
rect 2054 540 2071 557
rect 2054 506 2071 523
rect 2054 472 2071 489
rect 2054 438 2071 455
rect 2054 404 2071 421
rect 2054 370 2071 387
rect 2054 336 2071 353
rect 2054 302 2071 319
rect 2054 268 2071 285
rect 2054 234 2071 251
rect 2054 200 2071 217
rect 2054 166 2071 183
rect 2098 1118 2115 1135
rect 2098 1084 2115 1101
rect 2098 1050 2115 1067
rect 2098 1016 2115 1033
rect 2099 982 2116 999
rect 2099 948 2116 965
rect 2099 914 2116 931
rect 2099 880 2116 897
rect 2099 846 2116 863
rect 2099 812 2116 829
rect 2099 778 2116 795
rect 2099 744 2116 761
rect 2099 710 2116 727
rect 2099 676 2116 693
rect 2099 642 2116 659
rect 2099 608 2116 625
rect 2099 574 2116 591
rect 2099 540 2116 557
rect 2099 506 2116 523
rect 2099 472 2116 489
rect 2099 438 2116 455
rect 2099 404 2116 421
rect 2099 370 2116 387
rect 2099 336 2116 353
rect 2099 302 2116 319
rect 2099 268 2116 285
rect 2099 234 2116 251
rect 2099 200 2116 217
rect 2099 166 2116 183
rect 2143 1120 2160 1137
rect 2143 1086 2160 1103
rect 2143 1052 2160 1069
rect 2143 1018 2160 1035
rect 2143 984 2160 1001
rect 2143 950 2160 967
rect 2143 916 2160 933
rect 2143 882 2160 899
rect 2143 848 2160 865
rect 2143 814 2160 831
rect 2143 780 2160 797
rect 2143 746 2160 763
rect 2143 712 2160 729
rect 2143 678 2160 695
rect 2143 644 2160 661
rect 2143 610 2160 627
rect 2143 576 2160 593
rect 2143 542 2160 559
rect 2143 508 2160 525
rect 2143 474 2160 491
rect 2143 440 2160 457
rect 2143 406 2160 423
rect 2143 372 2160 389
rect 2143 338 2160 355
rect 2143 304 2160 321
rect 2143 270 2160 287
rect 2143 236 2160 253
rect 2143 202 2160 219
rect 2143 168 2160 185
rect 2187 1118 2204 1135
rect 2187 1084 2204 1101
rect 2187 1050 2204 1067
rect 2187 1016 2204 1033
rect 2188 982 2205 999
rect 2188 948 2205 965
rect 2188 914 2205 931
rect 2188 880 2205 897
rect 2188 846 2205 863
rect 2188 812 2205 829
rect 2188 778 2205 795
rect 2188 744 2205 761
rect 2188 710 2205 727
rect 2188 676 2205 693
rect 2188 642 2205 659
rect 2188 608 2205 625
rect 2188 574 2205 591
rect 2188 540 2205 557
rect 2188 506 2205 523
rect 2188 472 2205 489
rect 2188 438 2205 455
rect 2188 404 2205 421
rect 2188 370 2205 387
rect 2188 336 2205 353
rect 2188 302 2205 319
rect 2188 268 2205 285
rect 2188 234 2205 251
rect 2188 200 2205 217
rect 2188 166 2205 183
rect 2232 1118 2249 1135
rect 2232 1084 2249 1101
rect 2232 1050 2249 1067
rect 2232 1016 2249 1033
rect 2233 982 2250 999
rect 2233 948 2250 965
rect 2233 914 2250 931
rect 2233 880 2250 897
rect 2233 846 2250 863
rect 2233 812 2250 829
rect 2233 778 2250 795
rect 2233 744 2250 761
rect 2233 710 2250 727
rect 2233 676 2250 693
rect 2233 642 2250 659
rect 2233 608 2250 625
rect 2233 574 2250 591
rect 2233 540 2250 557
rect 2233 506 2250 523
rect 2233 472 2250 489
rect 2233 438 2250 455
rect 2233 404 2250 421
rect 2233 370 2250 387
rect 2233 336 2250 353
rect 2233 302 2250 319
rect 2233 268 2250 285
rect 2233 234 2250 251
rect 2233 200 2250 217
rect 2233 166 2250 183
rect 2277 1118 2294 1135
rect 2277 1084 2294 1101
rect 2277 1050 2294 1067
rect 2277 1016 2294 1033
rect 2278 982 2295 999
rect 2278 948 2295 965
rect 2278 914 2295 931
rect 2278 880 2295 897
rect 2278 846 2295 863
rect 2278 812 2295 829
rect 2278 778 2295 795
rect 2278 744 2295 761
rect 2278 710 2295 727
rect 2278 676 2295 693
rect 2278 642 2295 659
rect 2278 608 2295 625
rect 2278 574 2295 591
rect 2278 540 2295 557
rect 2278 506 2295 523
rect 2278 472 2295 489
rect 2278 438 2295 455
rect 2278 404 2295 421
rect 2278 370 2295 387
rect 2278 336 2295 353
rect 2278 302 2295 319
rect 2278 268 2295 285
rect 2278 234 2295 251
rect 2278 200 2295 217
rect 2278 166 2295 183
rect 2322 1118 2339 1135
rect 2322 1084 2339 1101
rect 2322 1050 2339 1067
rect 2322 1016 2339 1033
rect 2323 982 2340 999
rect 2323 948 2340 965
rect 2323 914 2340 931
rect 2323 880 2340 897
rect 2323 846 2340 863
rect 2323 812 2340 829
rect 2323 778 2340 795
rect 2323 744 2340 761
rect 2323 710 2340 727
rect 2323 676 2340 693
rect 2323 642 2340 659
rect 2323 608 2340 625
rect 2323 574 2340 591
rect 2323 540 2340 557
rect 2323 506 2340 523
rect 2323 472 2340 489
rect 2323 438 2340 455
rect 2323 404 2340 421
rect 2323 370 2340 387
rect 2323 336 2340 353
rect 2323 302 2340 319
rect 2323 268 2340 285
rect 2323 234 2340 251
rect 2323 200 2340 217
rect 2323 166 2340 183
rect 2367 1118 2384 1135
rect 2367 1084 2384 1101
rect 2367 1050 2384 1067
rect 2367 1016 2384 1033
rect 2368 982 2385 999
rect 2368 948 2385 965
rect 2368 914 2385 931
rect 2368 880 2385 897
rect 2368 846 2385 863
rect 2368 812 2385 829
rect 2368 778 2385 795
rect 2368 744 2385 761
rect 2368 710 2385 727
rect 2368 676 2385 693
rect 2368 642 2385 659
rect 2368 608 2385 625
rect 2368 574 2385 591
rect 2368 540 2385 557
rect 2368 506 2385 523
rect 2368 472 2385 489
rect 2368 438 2385 455
rect 2368 404 2385 421
rect 2368 370 2385 387
rect 2368 336 2385 353
rect 2368 302 2385 319
rect 2368 268 2385 285
rect 2368 234 2385 251
rect 2368 200 2385 217
rect 2368 166 2385 183
rect 2412 1118 2429 1135
rect 2412 1084 2429 1101
rect 2412 1050 2429 1067
rect 2412 1016 2429 1033
rect 2413 982 2430 999
rect 2413 948 2430 965
rect 2413 914 2430 931
rect 2413 880 2430 897
rect 2413 846 2430 863
rect 2413 812 2430 829
rect 2413 778 2430 795
rect 2413 744 2430 761
rect 2413 710 2430 727
rect 2413 676 2430 693
rect 2413 642 2430 659
rect 2413 608 2430 625
rect 2413 574 2430 591
rect 2413 540 2430 557
rect 2413 506 2430 523
rect 2413 472 2430 489
rect 2413 438 2430 455
rect 2413 404 2430 421
rect 2413 370 2430 387
rect 2413 336 2430 353
rect 2413 302 2430 319
rect 2413 268 2430 285
rect 2413 234 2430 251
rect 2413 200 2430 217
rect 2413 166 2430 183
rect 2458 1118 2475 1135
rect 2458 1084 2475 1101
rect 2458 1050 2475 1067
rect 2458 1016 2475 1033
rect 2459 982 2476 999
rect 2459 948 2476 965
rect 2459 914 2476 931
rect 2459 880 2476 897
rect 2459 846 2476 863
rect 2459 812 2476 829
rect 2459 778 2476 795
rect 2459 744 2476 761
rect 2459 710 2476 727
rect 2459 676 2476 693
rect 2459 642 2476 659
rect 2459 608 2476 625
rect 2459 574 2476 591
rect 2459 540 2476 557
rect 2459 506 2476 523
rect 2459 472 2476 489
rect 2459 438 2476 455
rect 2459 404 2476 421
rect 2459 370 2476 387
rect 2459 336 2476 353
rect 2459 302 2476 319
rect 2459 268 2476 285
rect 2459 234 2476 251
rect 2459 200 2476 217
rect 2459 166 2476 183
rect 2503 1120 2520 1137
rect 2503 1086 2520 1103
rect 2503 1052 2520 1069
rect 2503 1018 2520 1035
rect 2503 984 2520 1001
rect 2503 950 2520 967
rect 2503 916 2520 933
rect 2503 882 2520 899
rect 2503 848 2520 865
rect 2503 814 2520 831
rect 2503 780 2520 797
rect 2503 746 2520 763
rect 2503 712 2520 729
rect 2503 678 2520 695
rect 2503 644 2520 661
rect 2503 610 2520 627
rect 2503 576 2520 593
rect 2503 542 2520 559
rect 2503 508 2520 525
rect 2503 474 2520 491
rect 2503 440 2520 457
rect 2503 406 2520 423
rect 2503 372 2520 389
rect 2503 338 2520 355
rect 2503 304 2520 321
rect 2503 270 2520 287
rect 2503 236 2520 253
rect 2503 202 2520 219
rect 2503 168 2520 185
rect 2547 1118 2564 1135
rect 2547 1084 2564 1101
rect 2547 1050 2564 1067
rect 2547 1016 2564 1033
rect 2548 982 2565 999
rect 2548 948 2565 965
rect 2548 914 2565 931
rect 2548 880 2565 897
rect 2548 846 2565 863
rect 2548 812 2565 829
rect 2548 778 2565 795
rect 2548 744 2565 761
rect 2548 710 2565 727
rect 2548 676 2565 693
rect 2548 642 2565 659
rect 2548 608 2565 625
rect 2548 574 2565 591
rect 2548 540 2565 557
rect 2548 506 2565 523
rect 2548 472 2565 489
rect 2548 438 2565 455
rect 2548 404 2565 421
rect 2548 370 2565 387
rect 2548 336 2565 353
rect 2548 302 2565 319
rect 2548 268 2565 285
rect 2548 234 2565 251
rect 2548 200 2565 217
rect 2548 166 2565 183
rect 2592 1118 2609 1135
rect 2592 1084 2609 1101
rect 2592 1050 2609 1067
rect 2592 1016 2609 1033
rect 2593 982 2610 999
rect 2593 948 2610 965
rect 2593 914 2610 931
rect 2593 880 2610 897
rect 2593 846 2610 863
rect 2593 812 2610 829
rect 2593 778 2610 795
rect 2593 744 2610 761
rect 2593 710 2610 727
rect 2593 676 2610 693
rect 2593 642 2610 659
rect 2593 608 2610 625
rect 2593 574 2610 591
rect 2593 540 2610 557
rect 2593 506 2610 523
rect 2593 472 2610 489
rect 2593 438 2610 455
rect 2593 404 2610 421
rect 2593 370 2610 387
rect 2593 336 2610 353
rect 2593 302 2610 319
rect 2593 268 2610 285
rect 2593 234 2610 251
rect 2593 200 2610 217
rect 2593 166 2610 183
rect 2637 1118 2654 1135
rect 2637 1084 2654 1101
rect 2637 1050 2654 1067
rect 2637 1016 2654 1033
rect 2638 982 2655 999
rect 2638 948 2655 965
rect 2638 914 2655 931
rect 2638 880 2655 897
rect 2638 846 2655 863
rect 2638 812 2655 829
rect 2638 778 2655 795
rect 2638 744 2655 761
rect 2638 710 2655 727
rect 2638 676 2655 693
rect 2638 642 2655 659
rect 2638 608 2655 625
rect 2638 574 2655 591
rect 2638 540 2655 557
rect 2638 506 2655 523
rect 2638 472 2655 489
rect 2638 438 2655 455
rect 2638 404 2655 421
rect 2638 370 2655 387
rect 2638 336 2655 353
rect 2638 302 2655 319
rect 2638 268 2655 285
rect 2638 234 2655 251
rect 2638 200 2655 217
rect 2638 166 2655 183
<< psubdiff >>
rect -21 112 2613 121
rect -21 111 983 112
rect -21 110 641 111
rect -21 93 -9 110
rect 8 109 196 110
rect 8 93 25 109
rect -21 92 25 93
rect 42 92 59 109
rect 76 108 128 109
rect 76 92 94 108
rect -21 91 94 92
rect 111 92 128 108
rect 145 92 162 109
rect 179 93 196 109
rect 213 93 230 110
rect 247 93 265 110
rect 282 93 299 110
rect 316 109 470 110
rect 316 108 367 109
rect 316 93 333 108
rect 179 92 333 93
rect 111 91 333 92
rect 350 92 367 108
rect 384 92 401 109
rect 418 92 436 109
rect 453 93 470 109
rect 487 93 504 110
rect 521 93 538 110
rect 555 93 572 110
rect 589 93 607 110
rect 624 94 641 110
rect 658 110 812 111
rect 658 94 675 110
rect 624 93 675 94
rect 692 93 709 110
rect 726 93 743 110
rect 760 93 778 110
rect 795 94 812 110
rect 829 94 846 111
rect 863 94 880 111
rect 897 94 914 111
rect 931 94 949 111
rect 966 95 983 111
rect 1000 111 1256 112
rect 1000 95 1017 111
rect 966 94 1017 95
rect 1034 94 1051 111
rect 1068 94 1085 111
rect 1102 94 1120 111
rect 1137 94 1154 111
rect 1171 94 1188 111
rect 1205 94 1222 111
rect 1239 95 1256 111
rect 1273 111 1325 112
rect 1273 95 1291 111
rect 1239 94 1291 95
rect 1308 95 1325 111
rect 1342 110 1393 112
rect 1342 95 1359 110
rect 1308 94 1359 95
rect 795 93 1359 94
rect 1376 95 1393 110
rect 1410 111 1804 112
rect 1410 95 1427 111
rect 1376 94 1427 95
rect 1444 94 1462 111
rect 1479 94 1496 111
rect 1513 110 1633 111
rect 1513 94 1530 110
rect 1376 93 1530 94
rect 1547 93 1564 110
rect 1581 93 1599 110
rect 1616 94 1633 110
rect 1650 94 1667 111
rect 1684 94 1701 111
rect 1718 94 1735 111
rect 1752 94 1770 111
rect 1787 95 1804 111
rect 1821 111 1872 112
rect 1821 95 1838 111
rect 1787 94 1838 95
rect 1855 95 1872 111
rect 1889 111 1941 112
rect 1889 95 1906 111
rect 1855 94 1906 95
rect 1923 95 1941 111
rect 1958 111 2284 112
rect 1958 95 1976 111
rect 1923 94 1976 95
rect 1993 110 2079 111
rect 1993 94 2010 110
rect 1616 93 2010 94
rect 2027 93 2044 110
rect 2061 94 2079 110
rect 2096 94 2113 111
rect 2130 94 2147 111
rect 2164 94 2181 111
rect 2198 94 2215 111
rect 2232 94 2250 111
rect 2267 95 2284 111
rect 2301 111 2352 112
rect 2301 95 2318 111
rect 2267 94 2318 95
rect 2335 95 2352 111
rect 2369 111 2421 112
rect 2369 95 2386 111
rect 2335 94 2386 95
rect 2403 95 2421 111
rect 2438 111 2613 112
rect 2438 95 2455 111
rect 2403 94 2455 95
rect 2472 94 2489 111
rect 2506 110 2613 111
rect 2506 94 2523 110
rect 2061 93 2523 94
rect 2540 93 2558 110
rect 2575 108 2613 110
rect 2575 93 2592 108
rect 453 92 2592 93
rect 350 91 2592 92
rect 2609 91 2613 108
rect -21 79 2613 91
<< psubdiffcont >>
rect -9 93 8 110
rect 25 92 42 109
rect 59 92 76 109
rect 94 91 111 108
rect 128 92 145 109
rect 162 92 179 109
rect 196 93 213 110
rect 230 93 247 110
rect 265 93 282 110
rect 299 93 316 110
rect 333 91 350 108
rect 367 92 384 109
rect 401 92 418 109
rect 436 92 453 109
rect 470 93 487 110
rect 504 93 521 110
rect 538 93 555 110
rect 572 93 589 110
rect 607 93 624 110
rect 641 94 658 111
rect 675 93 692 110
rect 709 93 726 110
rect 743 93 760 110
rect 778 93 795 110
rect 812 94 829 111
rect 846 94 863 111
rect 880 94 897 111
rect 914 94 931 111
rect 949 94 966 111
rect 983 95 1000 112
rect 1017 94 1034 111
rect 1051 94 1068 111
rect 1085 94 1102 111
rect 1120 94 1137 111
rect 1154 94 1171 111
rect 1188 94 1205 111
rect 1222 94 1239 111
rect 1256 95 1273 112
rect 1291 94 1308 111
rect 1325 95 1342 112
rect 1359 93 1376 110
rect 1393 95 1410 112
rect 1427 94 1444 111
rect 1462 94 1479 111
rect 1496 94 1513 111
rect 1530 93 1547 110
rect 1564 93 1581 110
rect 1599 93 1616 110
rect 1633 94 1650 111
rect 1667 94 1684 111
rect 1701 94 1718 111
rect 1735 94 1752 111
rect 1770 94 1787 111
rect 1804 95 1821 112
rect 1838 94 1855 111
rect 1872 95 1889 112
rect 1906 94 1923 111
rect 1941 95 1958 112
rect 1976 94 1993 111
rect 2010 93 2027 110
rect 2044 93 2061 110
rect 2079 94 2096 111
rect 2113 94 2130 111
rect 2147 94 2164 111
rect 2181 94 2198 111
rect 2215 94 2232 111
rect 2250 94 2267 111
rect 2284 95 2301 112
rect 2318 94 2335 111
rect 2352 95 2369 112
rect 2386 94 2403 111
rect 2421 95 2438 112
rect 2455 94 2472 111
rect 2489 94 2506 111
rect 2523 93 2540 110
rect 2558 93 2575 110
rect 2592 91 2609 108
<< poly >>
rect -35 1161 24 1176
rect -35 1150 -20 1161
rect 9 1150 24 1161
rect 54 1161 114 1176
rect 54 1150 69 1161
rect 99 1150 114 1161
rect 144 1161 204 1176
rect 144 1150 159 1161
rect 189 1150 204 1161
rect 234 1161 294 1176
rect 234 1150 249 1161
rect 279 1150 294 1161
rect 325 1161 384 1176
rect 325 1150 340 1161
rect 369 1150 384 1161
rect 414 1161 474 1176
rect 414 1150 429 1161
rect 459 1150 474 1161
rect 504 1161 564 1176
rect 504 1150 519 1161
rect 549 1150 564 1161
rect 594 1161 654 1176
rect 594 1150 609 1161
rect 639 1150 654 1161
rect 684 1161 743 1176
rect 684 1150 699 1161
rect 728 1150 743 1161
rect 773 1161 833 1176
rect 773 1150 788 1161
rect 818 1150 833 1161
rect 863 1161 923 1176
rect 863 1150 878 1161
rect 908 1150 923 1161
rect 953 1161 1013 1176
rect 953 1150 968 1161
rect 998 1150 1013 1161
rect 1044 1161 1103 1176
rect 1044 1150 1059 1161
rect 1088 1150 1103 1161
rect 1133 1161 1193 1176
rect 1133 1150 1148 1161
rect 1178 1150 1193 1161
rect 1223 1161 1283 1176
rect 1223 1150 1238 1161
rect 1268 1150 1283 1161
rect 1313 1161 1373 1176
rect 1313 1150 1328 1161
rect 1358 1150 1373 1161
rect 1403 1161 1462 1176
rect 1403 1150 1418 1161
rect 1447 1150 1462 1161
rect 1492 1161 1552 1176
rect 1492 1150 1507 1161
rect 1537 1150 1552 1161
rect 1582 1161 1642 1176
rect 1582 1150 1597 1161
rect 1627 1150 1642 1161
rect 1672 1161 1732 1176
rect 1672 1150 1687 1161
rect 1717 1150 1732 1161
rect 1763 1161 1822 1176
rect 1763 1150 1778 1161
rect 1807 1150 1822 1161
rect 1852 1161 1912 1176
rect 1852 1150 1867 1161
rect 1897 1150 1912 1161
rect 1942 1161 2002 1176
rect 1942 1150 1957 1161
rect 1987 1150 2002 1161
rect 2032 1161 2092 1176
rect 2032 1150 2047 1161
rect 2077 1150 2092 1161
rect 2122 1161 2181 1176
rect 2122 1150 2137 1161
rect 2166 1150 2181 1161
rect 2211 1161 2271 1176
rect 2211 1150 2226 1161
rect 2256 1150 2271 1161
rect 2301 1161 2361 1176
rect 2301 1150 2316 1161
rect 2346 1150 2361 1161
rect 2391 1161 2451 1176
rect 2391 1150 2406 1161
rect 2436 1150 2451 1161
rect 2482 1161 2541 1176
rect 2482 1150 2497 1161
rect 2526 1150 2541 1161
rect 2571 1161 2631 1176
rect 2571 1150 2586 1161
rect 2616 1150 2631 1161
rect -196 142 -161 150
rect -35 142 -20 150
rect 9 142 24 150
rect 54 142 69 150
rect 99 142 114 150
rect 144 142 159 150
rect 189 142 204 150
rect 234 142 249 150
rect 279 142 294 150
rect 325 142 340 150
rect 369 142 384 150
rect 414 142 429 150
rect 459 142 474 150
rect 504 142 519 150
rect 549 142 564 150
rect 594 142 609 150
rect 639 142 654 150
rect 684 142 699 150
rect 728 142 743 150
rect 773 142 788 150
rect 818 142 833 150
rect 863 142 878 150
rect 908 142 923 150
rect 953 142 968 150
rect 998 142 1013 150
rect 1044 142 1059 150
rect 1088 142 1103 150
rect 1133 142 1148 150
rect 1178 142 1193 150
rect 1223 142 1238 150
rect 1268 142 1283 150
rect 1313 142 1328 150
rect 1358 142 1373 150
rect 1403 142 1418 150
rect 1447 142 1462 150
rect 1492 142 1507 150
rect 1537 142 1552 150
rect 1582 142 1597 150
rect 1627 142 1642 150
rect 1672 142 1687 150
rect 1717 142 1732 150
rect 1763 142 1778 150
rect 1807 142 1822 150
rect 1852 142 1867 150
rect 1897 142 1912 150
rect 1942 142 1957 150
rect 1987 142 2002 150
rect 2032 142 2047 150
rect 2077 142 2092 150
rect 2122 142 2137 150
rect 2166 142 2181 150
rect 2211 142 2226 150
rect 2256 142 2271 150
rect 2301 142 2316 150
rect 2346 142 2361 150
rect 2391 142 2406 150
rect 2436 142 2451 150
rect 2482 142 2497 150
rect 2526 142 2541 150
rect 2571 142 2586 150
rect 2616 142 2631 150
rect -196 141 2631 142
rect -196 122 -188 141
rect -168 127 2631 141
rect -168 122 -161 127
rect -196 114 -161 122
<< polycont >>
rect -188 122 -168 141
<< locali >>
rect -85 1220 2677 1253
rect -85 1203 -79 1220
rect -62 1203 -43 1220
rect -26 1219 2677 1220
rect -26 1203 -7 1219
rect -85 1202 -7 1203
rect 10 1202 29 1219
rect 46 1202 65 1219
rect 82 1202 101 1219
rect 118 1202 137 1219
rect 154 1202 173 1219
rect 190 1218 1185 1219
rect 190 1202 209 1218
rect -85 1201 209 1202
rect 226 1201 245 1218
rect 262 1201 281 1218
rect 298 1201 317 1218
rect 334 1201 354 1218
rect 371 1201 390 1218
rect 407 1217 787 1218
rect 407 1201 426 1217
rect -85 1200 426 1201
rect 443 1200 462 1217
rect 479 1200 498 1217
rect 515 1200 534 1217
rect 551 1200 570 1217
rect 587 1200 606 1217
rect 623 1216 787 1217
rect 623 1200 642 1216
rect -85 1199 642 1200
rect 659 1199 678 1216
rect 695 1199 714 1216
rect 731 1199 750 1216
rect 767 1201 787 1216
rect 804 1201 823 1218
rect 840 1201 859 1218
rect 876 1201 896 1218
rect 913 1201 932 1218
rect 949 1217 1185 1218
rect 949 1201 968 1217
rect 767 1200 968 1201
rect 985 1200 1004 1217
rect 1021 1200 1040 1217
rect 1057 1200 1076 1217
rect 1093 1200 1112 1217
rect 1129 1200 1148 1217
rect 1165 1202 1185 1217
rect 1202 1202 1221 1219
rect 1238 1202 1257 1219
rect 1274 1202 1294 1219
rect 1311 1202 1330 1219
rect 1347 1218 1582 1219
rect 1347 1202 1366 1218
rect 1165 1201 1366 1202
rect 1383 1201 1402 1218
rect 1419 1201 1438 1218
rect 1455 1201 1474 1218
rect 1491 1201 1510 1218
rect 1527 1201 1546 1218
rect 1563 1202 1582 1218
rect 1599 1202 1618 1219
rect 1635 1202 1654 1219
rect 1671 1202 1691 1219
rect 1708 1202 1727 1219
rect 1744 1218 1979 1219
rect 1744 1202 1763 1218
rect 1563 1201 1763 1202
rect 1780 1201 1799 1218
rect 1816 1201 1835 1218
rect 1852 1201 1871 1218
rect 1888 1201 1907 1218
rect 1924 1201 1943 1218
rect 1960 1202 1979 1218
rect 1996 1202 2015 1219
rect 2032 1202 2051 1219
rect 2068 1202 2088 1219
rect 2105 1202 2124 1219
rect 2141 1218 2376 1219
rect 2141 1202 2160 1218
rect 1960 1201 2160 1202
rect 2177 1201 2196 1218
rect 2213 1201 2232 1218
rect 2249 1201 2268 1218
rect 2285 1201 2304 1218
rect 2321 1201 2340 1218
rect 2357 1202 2376 1218
rect 2393 1202 2412 1219
rect 2429 1218 2677 1219
rect 2429 1202 2448 1218
rect 2357 1201 2448 1202
rect 2465 1201 2484 1218
rect 2501 1201 2525 1218
rect 2542 1201 2561 1218
rect 2578 1201 2601 1218
rect 2618 1201 2642 1218
rect 2659 1201 2677 1218
rect 1165 1200 2677 1201
rect 767 1199 2677 1200
rect -85 1195 2677 1199
rect -85 1194 2660 1195
rect -64 1184 2660 1194
rect -64 1135 -38 1184
rect -64 1118 -59 1135
rect -42 1118 -38 1135
rect -64 1101 -38 1118
rect -64 1084 -59 1101
rect -42 1084 -38 1101
rect -64 1067 -38 1084
rect -64 1050 -59 1067
rect -42 1050 -38 1067
rect -64 1033 -38 1050
rect -64 1016 -59 1033
rect -42 1016 -38 1033
rect -64 999 -38 1016
rect -64 982 -58 999
rect -41 982 -38 999
rect -64 965 -38 982
rect -64 948 -58 965
rect -41 948 -38 965
rect -64 931 -38 948
rect -64 914 -58 931
rect -41 914 -38 931
rect -64 897 -38 914
rect -64 880 -58 897
rect -41 880 -38 897
rect -64 863 -38 880
rect -64 846 -58 863
rect -41 846 -38 863
rect -64 829 -38 846
rect -64 812 -58 829
rect -41 812 -38 829
rect -64 795 -38 812
rect -64 778 -58 795
rect -41 778 -38 795
rect -64 761 -38 778
rect -64 744 -58 761
rect -41 744 -38 761
rect -64 727 -38 744
rect -64 710 -58 727
rect -41 710 -38 727
rect -64 693 -38 710
rect -64 676 -58 693
rect -41 676 -38 693
rect -64 659 -38 676
rect -64 642 -58 659
rect -41 642 -38 659
rect -64 625 -38 642
rect -64 608 -58 625
rect -41 608 -38 625
rect -64 591 -38 608
rect -64 574 -58 591
rect -41 574 -38 591
rect -64 557 -38 574
rect -64 540 -58 557
rect -41 540 -38 557
rect -64 523 -38 540
rect -64 506 -58 523
rect -41 506 -38 523
rect -64 489 -38 506
rect -64 472 -58 489
rect -41 472 -38 489
rect -64 455 -38 472
rect -64 438 -58 455
rect -41 438 -38 455
rect -64 421 -38 438
rect -64 404 -58 421
rect -41 404 -38 421
rect -64 387 -38 404
rect -64 370 -58 387
rect -41 370 -38 387
rect -64 353 -38 370
rect -64 336 -58 353
rect -41 336 -38 353
rect -64 319 -38 336
rect -64 302 -58 319
rect -41 302 -38 319
rect -64 285 -38 302
rect -64 268 -58 285
rect -41 268 -38 285
rect -64 251 -38 268
rect -64 234 -58 251
rect -41 234 -38 251
rect -64 217 -38 234
rect -64 200 -58 217
rect -41 200 -38 217
rect -64 183 -38 200
rect -64 166 -58 183
rect -41 166 -38 183
rect -64 158 -38 166
rect -17 1137 6 1145
rect -17 1120 -14 1137
rect 3 1120 6 1137
rect -17 1103 6 1120
rect -17 1086 -14 1103
rect 3 1086 6 1103
rect -17 1069 6 1086
rect -17 1052 -14 1069
rect 3 1052 6 1069
rect -17 1035 6 1052
rect -17 1018 -14 1035
rect 3 1018 6 1035
rect -17 1001 6 1018
rect -17 984 -14 1001
rect 3 984 6 1001
rect -17 967 6 984
rect -17 950 -14 967
rect 3 950 6 967
rect -17 933 6 950
rect -17 916 -14 933
rect 3 916 6 933
rect -17 899 6 916
rect -17 882 -14 899
rect 3 882 6 899
rect -17 865 6 882
rect -17 848 -14 865
rect 3 848 6 865
rect -17 831 6 848
rect -17 814 -14 831
rect 3 814 6 831
rect -17 797 6 814
rect -17 780 -14 797
rect 3 780 6 797
rect -17 763 6 780
rect -17 746 -14 763
rect 3 746 6 763
rect -17 729 6 746
rect -17 712 -14 729
rect 3 712 6 729
rect -17 695 6 712
rect -17 678 -14 695
rect 3 678 6 695
rect -17 661 6 678
rect -17 644 -14 661
rect 3 644 6 661
rect -17 627 6 644
rect -17 610 -14 627
rect 3 610 6 627
rect -17 593 6 610
rect -17 576 -14 593
rect 3 576 6 593
rect -17 559 6 576
rect -17 542 -14 559
rect 3 542 6 559
rect -17 525 6 542
rect -17 508 -14 525
rect 3 508 6 525
rect -17 491 6 508
rect -17 474 -14 491
rect 3 474 6 491
rect -17 457 6 474
rect -17 440 -14 457
rect 3 440 6 457
rect -17 423 6 440
rect -17 406 -14 423
rect 3 406 6 423
rect -17 389 6 406
rect -17 372 -14 389
rect 3 372 6 389
rect -17 355 6 372
rect -17 338 -14 355
rect 3 338 6 355
rect -17 321 6 338
rect -17 304 -14 321
rect 3 304 6 321
rect -17 287 6 304
rect -17 270 -14 287
rect 3 270 6 287
rect -17 253 6 270
rect -17 236 -14 253
rect 3 236 6 253
rect -17 219 6 236
rect -17 202 -14 219
rect 3 202 6 219
rect -17 185 6 202
rect -17 168 -14 185
rect 3 168 6 185
rect -260 141 -161 150
rect -260 123 -188 141
rect -196 122 -188 123
rect -168 122 -161 141
rect -196 114 -161 122
rect -17 115 6 168
rect 27 1135 51 1184
rect 27 1118 30 1135
rect 47 1118 51 1135
rect 27 1101 51 1118
rect 27 1084 30 1101
rect 47 1084 51 1101
rect 27 1067 51 1084
rect 27 1050 30 1067
rect 47 1050 51 1067
rect 27 1033 51 1050
rect 27 1016 30 1033
rect 47 1016 51 1033
rect 27 999 51 1016
rect 27 982 31 999
rect 48 982 51 999
rect 27 965 51 982
rect 27 948 31 965
rect 48 948 51 965
rect 27 931 51 948
rect 27 914 31 931
rect 48 914 51 931
rect 27 897 51 914
rect 27 880 31 897
rect 48 880 51 897
rect 27 863 51 880
rect 27 846 31 863
rect 48 846 51 863
rect 27 829 51 846
rect 27 812 31 829
rect 48 812 51 829
rect 27 795 51 812
rect 27 778 31 795
rect 48 778 51 795
rect 27 761 51 778
rect 27 744 31 761
rect 48 744 51 761
rect 27 727 51 744
rect 27 710 31 727
rect 48 710 51 727
rect 27 693 51 710
rect 27 676 31 693
rect 48 676 51 693
rect 27 659 51 676
rect 27 642 31 659
rect 48 642 51 659
rect 27 625 51 642
rect 27 608 31 625
rect 48 608 51 625
rect 27 591 51 608
rect 27 574 31 591
rect 48 574 51 591
rect 27 557 51 574
rect 27 540 31 557
rect 48 540 51 557
rect 27 523 51 540
rect 27 506 31 523
rect 48 506 51 523
rect 27 489 51 506
rect 27 472 31 489
rect 48 472 51 489
rect 27 455 51 472
rect 27 438 31 455
rect 48 438 51 455
rect 27 421 51 438
rect 27 404 31 421
rect 48 404 51 421
rect 27 387 51 404
rect 27 370 31 387
rect 48 370 51 387
rect 27 353 51 370
rect 27 336 31 353
rect 48 336 51 353
rect 27 319 51 336
rect 27 302 31 319
rect 48 302 51 319
rect 27 285 51 302
rect 27 268 31 285
rect 48 268 51 285
rect 27 251 51 268
rect 27 234 31 251
rect 48 234 51 251
rect 27 217 51 234
rect 27 200 31 217
rect 48 200 51 217
rect 27 183 51 200
rect 27 166 31 183
rect 48 166 51 183
rect 27 158 51 166
rect 72 1135 96 1143
rect 72 1118 75 1135
rect 92 1118 96 1135
rect 72 1101 96 1118
rect 72 1084 75 1101
rect 92 1084 96 1101
rect 72 1067 96 1084
rect 72 1050 75 1067
rect 92 1050 96 1067
rect 72 1033 96 1050
rect 72 1016 75 1033
rect 92 1016 96 1033
rect 72 999 96 1016
rect 72 982 76 999
rect 93 982 96 999
rect 72 965 96 982
rect 72 948 76 965
rect 93 948 96 965
rect 72 931 96 948
rect 72 914 76 931
rect 93 914 96 931
rect 72 897 96 914
rect 72 880 76 897
rect 93 880 96 897
rect 72 863 96 880
rect 72 846 76 863
rect 93 846 96 863
rect 72 829 96 846
rect 72 812 76 829
rect 93 812 96 829
rect 72 795 96 812
rect 72 778 76 795
rect 93 778 96 795
rect 72 761 96 778
rect 72 744 76 761
rect 93 744 96 761
rect 72 727 96 744
rect 72 710 76 727
rect 93 710 96 727
rect 72 693 96 710
rect 72 676 76 693
rect 93 676 96 693
rect 72 659 96 676
rect 72 642 76 659
rect 93 642 96 659
rect 72 625 96 642
rect 72 608 76 625
rect 93 608 96 625
rect 72 591 96 608
rect 72 574 76 591
rect 93 574 96 591
rect 72 557 96 574
rect 72 540 76 557
rect 93 540 96 557
rect 72 523 96 540
rect 72 506 76 523
rect 93 506 96 523
rect 72 489 96 506
rect 72 472 76 489
rect 93 472 96 489
rect 72 455 96 472
rect 72 438 76 455
rect 93 438 96 455
rect 72 421 96 438
rect 72 404 76 421
rect 93 404 96 421
rect 72 387 96 404
rect 72 370 76 387
rect 93 370 96 387
rect 72 353 96 370
rect 72 336 76 353
rect 93 336 96 353
rect 72 319 96 336
rect 72 302 76 319
rect 93 302 96 319
rect 72 285 96 302
rect 72 268 76 285
rect 93 268 96 285
rect 72 251 96 268
rect 72 234 76 251
rect 93 234 96 251
rect 72 217 96 234
rect 72 200 76 217
rect 93 200 96 217
rect 72 183 96 200
rect 72 166 76 183
rect 93 166 96 183
rect 72 115 96 166
rect 117 1135 141 1184
rect 117 1118 120 1135
rect 137 1118 141 1135
rect 117 1101 141 1118
rect 117 1084 120 1101
rect 137 1084 141 1101
rect 117 1067 141 1084
rect 117 1050 120 1067
rect 137 1050 141 1067
rect 117 1033 141 1050
rect 117 1016 120 1033
rect 137 1016 141 1033
rect 117 999 141 1016
rect 117 982 121 999
rect 138 982 141 999
rect 117 965 141 982
rect 117 948 121 965
rect 138 948 141 965
rect 117 931 141 948
rect 117 914 121 931
rect 138 914 141 931
rect 117 897 141 914
rect 117 880 121 897
rect 138 880 141 897
rect 117 863 141 880
rect 117 846 121 863
rect 138 846 141 863
rect 117 829 141 846
rect 117 812 121 829
rect 138 812 141 829
rect 117 795 141 812
rect 117 778 121 795
rect 138 778 141 795
rect 117 761 141 778
rect 117 744 121 761
rect 138 744 141 761
rect 117 727 141 744
rect 117 710 121 727
rect 138 710 141 727
rect 117 693 141 710
rect 117 676 121 693
rect 138 676 141 693
rect 117 659 141 676
rect 117 642 121 659
rect 138 642 141 659
rect 117 625 141 642
rect 117 608 121 625
rect 138 608 141 625
rect 117 591 141 608
rect 117 574 121 591
rect 138 574 141 591
rect 117 557 141 574
rect 117 540 121 557
rect 138 540 141 557
rect 117 523 141 540
rect 117 506 121 523
rect 138 506 141 523
rect 117 489 141 506
rect 117 472 121 489
rect 138 472 141 489
rect 117 455 141 472
rect 117 438 121 455
rect 138 438 141 455
rect 117 421 141 438
rect 117 404 121 421
rect 138 404 141 421
rect 117 387 141 404
rect 117 370 121 387
rect 138 370 141 387
rect 117 353 141 370
rect 117 336 121 353
rect 138 336 141 353
rect 117 319 141 336
rect 117 302 121 319
rect 138 302 141 319
rect 117 285 141 302
rect 117 268 121 285
rect 138 268 141 285
rect 117 251 141 268
rect 117 234 121 251
rect 138 234 141 251
rect 117 217 141 234
rect 117 200 121 217
rect 138 200 141 217
rect 117 183 141 200
rect 117 166 121 183
rect 138 166 141 183
rect 117 158 141 166
rect 162 1135 186 1143
rect 162 1118 165 1135
rect 182 1118 186 1135
rect 162 1101 186 1118
rect 162 1084 165 1101
rect 182 1084 186 1101
rect 162 1067 186 1084
rect 162 1050 165 1067
rect 182 1050 186 1067
rect 162 1033 186 1050
rect 162 1016 165 1033
rect 182 1016 186 1033
rect 162 999 186 1016
rect 162 982 166 999
rect 183 982 186 999
rect 162 965 186 982
rect 162 948 166 965
rect 183 948 186 965
rect 162 931 186 948
rect 162 914 166 931
rect 183 914 186 931
rect 162 897 186 914
rect 162 880 166 897
rect 183 880 186 897
rect 162 863 186 880
rect 162 846 166 863
rect 183 846 186 863
rect 162 829 186 846
rect 162 812 166 829
rect 183 812 186 829
rect 162 795 186 812
rect 162 778 166 795
rect 183 778 186 795
rect 162 761 186 778
rect 162 744 166 761
rect 183 744 186 761
rect 162 727 186 744
rect 162 710 166 727
rect 183 710 186 727
rect 162 693 186 710
rect 162 676 166 693
rect 183 676 186 693
rect 162 659 186 676
rect 162 642 166 659
rect 183 642 186 659
rect 162 625 186 642
rect 162 608 166 625
rect 183 608 186 625
rect 162 591 186 608
rect 162 574 166 591
rect 183 574 186 591
rect 162 557 186 574
rect 162 540 166 557
rect 183 540 186 557
rect 162 523 186 540
rect 162 506 166 523
rect 183 506 186 523
rect 162 489 186 506
rect 162 472 166 489
rect 183 472 186 489
rect 162 455 186 472
rect 162 438 166 455
rect 183 438 186 455
rect 162 421 186 438
rect 162 404 166 421
rect 183 404 186 421
rect 162 387 186 404
rect 162 370 166 387
rect 183 370 186 387
rect 162 353 186 370
rect 162 336 166 353
rect 183 336 186 353
rect 162 319 186 336
rect 162 302 166 319
rect 183 302 186 319
rect 162 285 186 302
rect 162 268 166 285
rect 183 268 186 285
rect 162 251 186 268
rect 162 234 166 251
rect 183 234 186 251
rect 162 217 186 234
rect 162 200 166 217
rect 183 200 186 217
rect 162 183 186 200
rect 162 166 166 183
rect 183 166 186 183
rect 162 115 186 166
rect 207 1135 231 1184
rect 207 1118 210 1135
rect 227 1118 231 1135
rect 207 1101 231 1118
rect 207 1084 210 1101
rect 227 1084 231 1101
rect 207 1067 231 1084
rect 207 1050 210 1067
rect 227 1050 231 1067
rect 207 1033 231 1050
rect 207 1016 210 1033
rect 227 1016 231 1033
rect 207 999 231 1016
rect 207 982 211 999
rect 228 982 231 999
rect 207 965 231 982
rect 207 948 211 965
rect 228 948 231 965
rect 207 931 231 948
rect 207 914 211 931
rect 228 914 231 931
rect 207 897 231 914
rect 207 880 211 897
rect 228 880 231 897
rect 207 863 231 880
rect 207 846 211 863
rect 228 846 231 863
rect 207 829 231 846
rect 207 812 211 829
rect 228 812 231 829
rect 207 795 231 812
rect 207 778 211 795
rect 228 778 231 795
rect 207 761 231 778
rect 207 744 211 761
rect 228 744 231 761
rect 207 727 231 744
rect 207 710 211 727
rect 228 710 231 727
rect 207 693 231 710
rect 207 676 211 693
rect 228 676 231 693
rect 207 659 231 676
rect 207 642 211 659
rect 228 642 231 659
rect 207 625 231 642
rect 207 608 211 625
rect 228 608 231 625
rect 207 591 231 608
rect 207 574 211 591
rect 228 574 231 591
rect 207 557 231 574
rect 207 540 211 557
rect 228 540 231 557
rect 207 523 231 540
rect 207 506 211 523
rect 228 506 231 523
rect 207 489 231 506
rect 207 472 211 489
rect 228 472 231 489
rect 207 455 231 472
rect 207 438 211 455
rect 228 438 231 455
rect 207 421 231 438
rect 207 404 211 421
rect 228 404 231 421
rect 207 387 231 404
rect 207 370 211 387
rect 228 370 231 387
rect 207 353 231 370
rect 207 336 211 353
rect 228 336 231 353
rect 207 319 231 336
rect 207 302 211 319
rect 228 302 231 319
rect 207 285 231 302
rect 207 268 211 285
rect 228 268 231 285
rect 207 251 231 268
rect 207 234 211 251
rect 228 234 231 251
rect 207 217 231 234
rect 207 200 211 217
rect 228 200 231 217
rect 207 183 231 200
rect 207 166 211 183
rect 228 166 231 183
rect 207 158 231 166
rect 252 1135 276 1143
rect 252 1118 255 1135
rect 272 1118 276 1135
rect 252 1101 276 1118
rect 252 1084 255 1101
rect 272 1084 276 1101
rect 252 1067 276 1084
rect 252 1050 255 1067
rect 272 1050 276 1067
rect 252 1033 276 1050
rect 252 1016 255 1033
rect 272 1016 276 1033
rect 252 999 276 1016
rect 252 982 256 999
rect 273 982 276 999
rect 252 965 276 982
rect 252 948 256 965
rect 273 948 276 965
rect 252 931 276 948
rect 252 914 256 931
rect 273 914 276 931
rect 252 897 276 914
rect 252 880 256 897
rect 273 880 276 897
rect 252 863 276 880
rect 252 846 256 863
rect 273 846 276 863
rect 252 829 276 846
rect 252 812 256 829
rect 273 812 276 829
rect 252 795 276 812
rect 252 778 256 795
rect 273 778 276 795
rect 252 761 276 778
rect 252 744 256 761
rect 273 744 276 761
rect 252 727 276 744
rect 252 710 256 727
rect 273 710 276 727
rect 252 693 276 710
rect 252 676 256 693
rect 273 676 276 693
rect 252 659 276 676
rect 252 642 256 659
rect 273 642 276 659
rect 252 625 276 642
rect 252 608 256 625
rect 273 608 276 625
rect 252 591 276 608
rect 252 574 256 591
rect 273 574 276 591
rect 252 557 276 574
rect 252 540 256 557
rect 273 540 276 557
rect 252 523 276 540
rect 252 506 256 523
rect 273 506 276 523
rect 252 489 276 506
rect 252 472 256 489
rect 273 472 276 489
rect 252 455 276 472
rect 252 438 256 455
rect 273 438 276 455
rect 252 421 276 438
rect 252 404 256 421
rect 273 404 276 421
rect 252 387 276 404
rect 252 370 256 387
rect 273 370 276 387
rect 252 353 276 370
rect 252 336 256 353
rect 273 336 276 353
rect 252 319 276 336
rect 252 302 256 319
rect 273 302 276 319
rect 252 285 276 302
rect 252 268 256 285
rect 273 268 276 285
rect 252 251 276 268
rect 252 234 256 251
rect 273 234 276 251
rect 252 217 276 234
rect 252 200 256 217
rect 273 200 276 217
rect 252 183 276 200
rect 252 166 256 183
rect 273 166 276 183
rect 252 115 276 166
rect 298 1135 322 1184
rect 298 1118 301 1135
rect 318 1118 322 1135
rect 298 1101 322 1118
rect 298 1084 301 1101
rect 318 1084 322 1101
rect 298 1067 322 1084
rect 298 1050 301 1067
rect 318 1050 322 1067
rect 298 1033 322 1050
rect 298 1016 301 1033
rect 318 1016 322 1033
rect 298 999 322 1016
rect 298 982 302 999
rect 319 982 322 999
rect 298 965 322 982
rect 298 948 302 965
rect 319 948 322 965
rect 298 931 322 948
rect 298 914 302 931
rect 319 914 322 931
rect 298 897 322 914
rect 298 880 302 897
rect 319 880 322 897
rect 298 863 322 880
rect 298 846 302 863
rect 319 846 322 863
rect 298 829 322 846
rect 298 812 302 829
rect 319 812 322 829
rect 298 795 322 812
rect 298 778 302 795
rect 319 778 322 795
rect 298 761 322 778
rect 298 744 302 761
rect 319 744 322 761
rect 298 727 322 744
rect 298 710 302 727
rect 319 710 322 727
rect 298 693 322 710
rect 298 676 302 693
rect 319 676 322 693
rect 298 659 322 676
rect 298 642 302 659
rect 319 642 322 659
rect 298 625 322 642
rect 298 608 302 625
rect 319 608 322 625
rect 298 591 322 608
rect 298 574 302 591
rect 319 574 322 591
rect 298 557 322 574
rect 298 540 302 557
rect 319 540 322 557
rect 298 523 322 540
rect 298 506 302 523
rect 319 506 322 523
rect 298 489 322 506
rect 298 472 302 489
rect 319 472 322 489
rect 298 455 322 472
rect 298 438 302 455
rect 319 438 322 455
rect 298 421 322 438
rect 298 404 302 421
rect 319 404 322 421
rect 298 387 322 404
rect 298 370 302 387
rect 319 370 322 387
rect 298 353 322 370
rect 298 336 302 353
rect 319 336 322 353
rect 298 319 322 336
rect 298 302 302 319
rect 319 302 322 319
rect 298 285 322 302
rect 298 268 302 285
rect 319 268 322 285
rect 298 251 322 268
rect 298 234 302 251
rect 319 234 322 251
rect 298 217 322 234
rect 298 200 302 217
rect 319 200 322 217
rect 298 183 322 200
rect 298 166 302 183
rect 319 166 322 183
rect 298 158 322 166
rect 343 1137 366 1145
rect 343 1120 346 1137
rect 363 1120 366 1137
rect 343 1103 366 1120
rect 343 1086 346 1103
rect 363 1086 366 1103
rect 343 1069 366 1086
rect 343 1052 346 1069
rect 363 1052 366 1069
rect 343 1035 366 1052
rect 343 1018 346 1035
rect 363 1018 366 1035
rect 343 1001 366 1018
rect 343 984 346 1001
rect 363 984 366 1001
rect 343 967 366 984
rect 343 950 346 967
rect 363 950 366 967
rect 343 933 366 950
rect 343 916 346 933
rect 363 916 366 933
rect 343 899 366 916
rect 343 882 346 899
rect 363 882 366 899
rect 343 865 366 882
rect 343 848 346 865
rect 363 848 366 865
rect 343 831 366 848
rect 343 814 346 831
rect 363 814 366 831
rect 343 797 366 814
rect 343 780 346 797
rect 363 780 366 797
rect 343 763 366 780
rect 343 746 346 763
rect 363 746 366 763
rect 343 729 366 746
rect 343 712 346 729
rect 363 712 366 729
rect 343 695 366 712
rect 343 678 346 695
rect 363 678 366 695
rect 343 661 366 678
rect 343 644 346 661
rect 363 644 366 661
rect 343 627 366 644
rect 343 610 346 627
rect 363 610 366 627
rect 343 593 366 610
rect 343 576 346 593
rect 363 576 366 593
rect 343 559 366 576
rect 343 542 346 559
rect 363 542 366 559
rect 343 525 366 542
rect 343 508 346 525
rect 363 508 366 525
rect 343 491 366 508
rect 343 474 346 491
rect 363 474 366 491
rect 343 457 366 474
rect 343 440 346 457
rect 363 440 366 457
rect 343 423 366 440
rect 343 406 346 423
rect 363 406 366 423
rect 343 389 366 406
rect 343 372 346 389
rect 363 372 366 389
rect 343 355 366 372
rect 343 338 346 355
rect 363 338 366 355
rect 343 321 366 338
rect 343 304 346 321
rect 363 304 366 321
rect 343 287 366 304
rect 343 270 346 287
rect 363 270 366 287
rect 343 253 366 270
rect 343 236 346 253
rect 363 236 366 253
rect 343 219 366 236
rect 343 202 346 219
rect 363 202 366 219
rect 343 185 366 202
rect 343 168 346 185
rect 363 168 366 185
rect 343 115 366 168
rect 387 1135 411 1184
rect 387 1118 390 1135
rect 407 1118 411 1135
rect 387 1101 411 1118
rect 387 1084 390 1101
rect 407 1084 411 1101
rect 387 1067 411 1084
rect 387 1050 390 1067
rect 407 1050 411 1067
rect 387 1033 411 1050
rect 387 1016 390 1033
rect 407 1016 411 1033
rect 387 999 411 1016
rect 387 982 391 999
rect 408 982 411 999
rect 387 965 411 982
rect 387 948 391 965
rect 408 948 411 965
rect 387 931 411 948
rect 387 914 391 931
rect 408 914 411 931
rect 387 897 411 914
rect 387 880 391 897
rect 408 880 411 897
rect 387 863 411 880
rect 387 846 391 863
rect 408 846 411 863
rect 387 829 411 846
rect 387 812 391 829
rect 408 812 411 829
rect 387 795 411 812
rect 387 778 391 795
rect 408 778 411 795
rect 387 761 411 778
rect 387 744 391 761
rect 408 744 411 761
rect 387 727 411 744
rect 387 710 391 727
rect 408 710 411 727
rect 387 693 411 710
rect 387 676 391 693
rect 408 676 411 693
rect 387 659 411 676
rect 387 642 391 659
rect 408 642 411 659
rect 387 625 411 642
rect 387 608 391 625
rect 408 608 411 625
rect 387 591 411 608
rect 387 574 391 591
rect 408 574 411 591
rect 387 557 411 574
rect 387 540 391 557
rect 408 540 411 557
rect 387 523 411 540
rect 387 506 391 523
rect 408 506 411 523
rect 387 489 411 506
rect 387 472 391 489
rect 408 472 411 489
rect 387 455 411 472
rect 387 438 391 455
rect 408 438 411 455
rect 387 421 411 438
rect 387 404 391 421
rect 408 404 411 421
rect 387 387 411 404
rect 387 370 391 387
rect 408 370 411 387
rect 387 353 411 370
rect 387 336 391 353
rect 408 336 411 353
rect 387 319 411 336
rect 387 302 391 319
rect 408 302 411 319
rect 387 285 411 302
rect 387 268 391 285
rect 408 268 411 285
rect 387 251 411 268
rect 387 234 391 251
rect 408 234 411 251
rect 387 217 411 234
rect 387 200 391 217
rect 408 200 411 217
rect 387 183 411 200
rect 387 166 391 183
rect 408 166 411 183
rect 387 158 411 166
rect 432 1135 456 1143
rect 432 1118 435 1135
rect 452 1118 456 1135
rect 432 1101 456 1118
rect 432 1084 435 1101
rect 452 1084 456 1101
rect 432 1067 456 1084
rect 432 1050 435 1067
rect 452 1050 456 1067
rect 432 1033 456 1050
rect 432 1016 435 1033
rect 452 1016 456 1033
rect 432 999 456 1016
rect 432 982 436 999
rect 453 982 456 999
rect 432 965 456 982
rect 432 948 436 965
rect 453 948 456 965
rect 432 931 456 948
rect 432 914 436 931
rect 453 914 456 931
rect 432 897 456 914
rect 432 880 436 897
rect 453 880 456 897
rect 432 863 456 880
rect 432 846 436 863
rect 453 846 456 863
rect 432 829 456 846
rect 432 812 436 829
rect 453 812 456 829
rect 432 795 456 812
rect 432 778 436 795
rect 453 778 456 795
rect 432 761 456 778
rect 432 744 436 761
rect 453 744 456 761
rect 432 727 456 744
rect 432 710 436 727
rect 453 710 456 727
rect 432 693 456 710
rect 432 676 436 693
rect 453 676 456 693
rect 432 659 456 676
rect 432 642 436 659
rect 453 642 456 659
rect 432 625 456 642
rect 432 608 436 625
rect 453 608 456 625
rect 432 591 456 608
rect 432 574 436 591
rect 453 574 456 591
rect 432 557 456 574
rect 432 540 436 557
rect 453 540 456 557
rect 432 523 456 540
rect 432 506 436 523
rect 453 506 456 523
rect 432 489 456 506
rect 432 472 436 489
rect 453 472 456 489
rect 432 455 456 472
rect 432 438 436 455
rect 453 438 456 455
rect 432 421 456 438
rect 432 404 436 421
rect 453 404 456 421
rect 432 387 456 404
rect 432 370 436 387
rect 453 370 456 387
rect 432 353 456 370
rect 432 336 436 353
rect 453 336 456 353
rect 432 319 456 336
rect 432 302 436 319
rect 453 302 456 319
rect 432 285 456 302
rect 432 268 436 285
rect 453 268 456 285
rect 432 251 456 268
rect 432 234 436 251
rect 453 234 456 251
rect 432 217 456 234
rect 432 200 436 217
rect 453 200 456 217
rect 432 183 456 200
rect 432 166 436 183
rect 453 166 456 183
rect 432 115 456 166
rect 477 1135 501 1184
rect 477 1118 480 1135
rect 497 1118 501 1135
rect 477 1101 501 1118
rect 477 1084 480 1101
rect 497 1084 501 1101
rect 477 1067 501 1084
rect 477 1050 480 1067
rect 497 1050 501 1067
rect 477 1033 501 1050
rect 477 1016 480 1033
rect 497 1016 501 1033
rect 477 999 501 1016
rect 477 982 481 999
rect 498 982 501 999
rect 477 965 501 982
rect 477 948 481 965
rect 498 948 501 965
rect 477 931 501 948
rect 477 914 481 931
rect 498 914 501 931
rect 477 897 501 914
rect 477 880 481 897
rect 498 880 501 897
rect 477 863 501 880
rect 477 846 481 863
rect 498 846 501 863
rect 477 829 501 846
rect 477 812 481 829
rect 498 812 501 829
rect 477 795 501 812
rect 477 778 481 795
rect 498 778 501 795
rect 477 761 501 778
rect 477 744 481 761
rect 498 744 501 761
rect 477 727 501 744
rect 477 710 481 727
rect 498 710 501 727
rect 477 693 501 710
rect 477 676 481 693
rect 498 676 501 693
rect 477 659 501 676
rect 477 642 481 659
rect 498 642 501 659
rect 477 625 501 642
rect 477 608 481 625
rect 498 608 501 625
rect 477 591 501 608
rect 477 574 481 591
rect 498 574 501 591
rect 477 557 501 574
rect 477 540 481 557
rect 498 540 501 557
rect 477 523 501 540
rect 477 506 481 523
rect 498 506 501 523
rect 477 489 501 506
rect 477 472 481 489
rect 498 472 501 489
rect 477 455 501 472
rect 477 438 481 455
rect 498 438 501 455
rect 477 421 501 438
rect 477 404 481 421
rect 498 404 501 421
rect 477 387 501 404
rect 477 370 481 387
rect 498 370 501 387
rect 477 353 501 370
rect 477 336 481 353
rect 498 336 501 353
rect 477 319 501 336
rect 477 302 481 319
rect 498 302 501 319
rect 477 285 501 302
rect 477 268 481 285
rect 498 268 501 285
rect 477 251 501 268
rect 477 234 481 251
rect 498 234 501 251
rect 477 217 501 234
rect 477 200 481 217
rect 498 200 501 217
rect 477 183 501 200
rect 477 166 481 183
rect 498 166 501 183
rect 477 158 501 166
rect 522 1135 546 1143
rect 522 1118 525 1135
rect 542 1118 546 1135
rect 522 1101 546 1118
rect 522 1084 525 1101
rect 542 1084 546 1101
rect 522 1067 546 1084
rect 522 1050 525 1067
rect 542 1050 546 1067
rect 522 1033 546 1050
rect 522 1016 525 1033
rect 542 1016 546 1033
rect 522 999 546 1016
rect 522 982 526 999
rect 543 982 546 999
rect 522 965 546 982
rect 522 948 526 965
rect 543 948 546 965
rect 522 931 546 948
rect 522 914 526 931
rect 543 914 546 931
rect 522 897 546 914
rect 522 880 526 897
rect 543 880 546 897
rect 522 863 546 880
rect 522 846 526 863
rect 543 846 546 863
rect 522 829 546 846
rect 522 812 526 829
rect 543 812 546 829
rect 522 795 546 812
rect 522 778 526 795
rect 543 778 546 795
rect 522 761 546 778
rect 522 744 526 761
rect 543 744 546 761
rect 522 727 546 744
rect 522 710 526 727
rect 543 710 546 727
rect 522 693 546 710
rect 522 676 526 693
rect 543 676 546 693
rect 522 659 546 676
rect 522 642 526 659
rect 543 642 546 659
rect 522 625 546 642
rect 522 608 526 625
rect 543 608 546 625
rect 522 591 546 608
rect 522 574 526 591
rect 543 574 546 591
rect 522 557 546 574
rect 522 540 526 557
rect 543 540 546 557
rect 522 523 546 540
rect 522 506 526 523
rect 543 506 546 523
rect 522 489 546 506
rect 522 472 526 489
rect 543 472 546 489
rect 522 455 546 472
rect 522 438 526 455
rect 543 438 546 455
rect 522 421 546 438
rect 522 404 526 421
rect 543 404 546 421
rect 522 387 546 404
rect 522 370 526 387
rect 543 370 546 387
rect 522 353 546 370
rect 522 336 526 353
rect 543 336 546 353
rect 522 319 546 336
rect 522 302 526 319
rect 543 302 546 319
rect 522 285 546 302
rect 522 268 526 285
rect 543 268 546 285
rect 522 251 546 268
rect 522 234 526 251
rect 543 234 546 251
rect 522 217 546 234
rect 522 200 526 217
rect 543 200 546 217
rect 522 183 546 200
rect 522 166 526 183
rect 543 166 546 183
rect 522 115 546 166
rect 567 1135 591 1184
rect 567 1118 570 1135
rect 587 1118 591 1135
rect 567 1101 591 1118
rect 567 1084 570 1101
rect 587 1084 591 1101
rect 567 1067 591 1084
rect 567 1050 570 1067
rect 587 1050 591 1067
rect 567 1033 591 1050
rect 567 1016 570 1033
rect 587 1016 591 1033
rect 567 999 591 1016
rect 567 982 571 999
rect 588 982 591 999
rect 567 965 591 982
rect 567 948 571 965
rect 588 948 591 965
rect 567 931 591 948
rect 567 914 571 931
rect 588 914 591 931
rect 567 897 591 914
rect 567 880 571 897
rect 588 880 591 897
rect 567 863 591 880
rect 567 846 571 863
rect 588 846 591 863
rect 567 829 591 846
rect 567 812 571 829
rect 588 812 591 829
rect 567 795 591 812
rect 567 778 571 795
rect 588 778 591 795
rect 567 761 591 778
rect 567 744 571 761
rect 588 744 591 761
rect 567 727 591 744
rect 567 710 571 727
rect 588 710 591 727
rect 567 693 591 710
rect 567 676 571 693
rect 588 676 591 693
rect 567 659 591 676
rect 567 642 571 659
rect 588 642 591 659
rect 567 625 591 642
rect 567 608 571 625
rect 588 608 591 625
rect 567 591 591 608
rect 567 574 571 591
rect 588 574 591 591
rect 567 557 591 574
rect 567 540 571 557
rect 588 540 591 557
rect 567 523 591 540
rect 567 506 571 523
rect 588 506 591 523
rect 567 489 591 506
rect 567 472 571 489
rect 588 472 591 489
rect 567 455 591 472
rect 567 438 571 455
rect 588 438 591 455
rect 567 421 591 438
rect 567 404 571 421
rect 588 404 591 421
rect 567 387 591 404
rect 567 370 571 387
rect 588 370 591 387
rect 567 353 591 370
rect 567 336 571 353
rect 588 336 591 353
rect 567 319 591 336
rect 567 302 571 319
rect 588 302 591 319
rect 567 285 591 302
rect 567 268 571 285
rect 588 268 591 285
rect 567 251 591 268
rect 567 234 571 251
rect 588 234 591 251
rect 567 217 591 234
rect 567 200 571 217
rect 588 200 591 217
rect 567 183 591 200
rect 567 166 571 183
rect 588 166 591 183
rect 567 158 591 166
rect 612 1135 636 1143
rect 612 1118 615 1135
rect 632 1118 636 1135
rect 612 1101 636 1118
rect 612 1084 615 1101
rect 632 1084 636 1101
rect 612 1067 636 1084
rect 612 1050 615 1067
rect 632 1050 636 1067
rect 612 1033 636 1050
rect 612 1016 615 1033
rect 632 1016 636 1033
rect 612 999 636 1016
rect 612 982 616 999
rect 633 982 636 999
rect 612 965 636 982
rect 612 948 616 965
rect 633 948 636 965
rect 612 931 636 948
rect 612 914 616 931
rect 633 914 636 931
rect 612 897 636 914
rect 612 880 616 897
rect 633 880 636 897
rect 612 863 636 880
rect 612 846 616 863
rect 633 846 636 863
rect 612 829 636 846
rect 612 812 616 829
rect 633 812 636 829
rect 612 795 636 812
rect 612 778 616 795
rect 633 778 636 795
rect 612 761 636 778
rect 612 744 616 761
rect 633 744 636 761
rect 612 727 636 744
rect 612 710 616 727
rect 633 710 636 727
rect 612 693 636 710
rect 612 676 616 693
rect 633 676 636 693
rect 612 659 636 676
rect 612 642 616 659
rect 633 642 636 659
rect 612 625 636 642
rect 612 608 616 625
rect 633 608 636 625
rect 612 591 636 608
rect 612 574 616 591
rect 633 574 636 591
rect 612 557 636 574
rect 612 540 616 557
rect 633 540 636 557
rect 612 523 636 540
rect 612 506 616 523
rect 633 506 636 523
rect 612 489 636 506
rect 612 472 616 489
rect 633 472 636 489
rect 612 455 636 472
rect 612 438 616 455
rect 633 438 636 455
rect 612 421 636 438
rect 612 404 616 421
rect 633 404 636 421
rect 612 387 636 404
rect 612 370 616 387
rect 633 370 636 387
rect 612 353 636 370
rect 612 336 616 353
rect 633 336 636 353
rect 612 319 636 336
rect 612 302 616 319
rect 633 302 636 319
rect 612 285 636 302
rect 612 268 616 285
rect 633 268 636 285
rect 612 251 636 268
rect 612 234 616 251
rect 633 234 636 251
rect 612 217 636 234
rect 612 200 616 217
rect 633 200 636 217
rect 612 183 636 200
rect 612 166 616 183
rect 633 166 636 183
rect 612 115 636 166
rect 657 1135 681 1184
rect 657 1118 660 1135
rect 677 1118 681 1135
rect 657 1101 681 1118
rect 657 1084 660 1101
rect 677 1084 681 1101
rect 657 1067 681 1084
rect 657 1050 660 1067
rect 677 1050 681 1067
rect 657 1033 681 1050
rect 657 1016 660 1033
rect 677 1016 681 1033
rect 657 999 681 1016
rect 657 982 661 999
rect 678 982 681 999
rect 657 965 681 982
rect 657 948 661 965
rect 678 948 681 965
rect 657 931 681 948
rect 657 914 661 931
rect 678 914 681 931
rect 657 897 681 914
rect 657 880 661 897
rect 678 880 681 897
rect 657 863 681 880
rect 657 846 661 863
rect 678 846 681 863
rect 657 829 681 846
rect 657 812 661 829
rect 678 812 681 829
rect 657 795 681 812
rect 657 778 661 795
rect 678 778 681 795
rect 657 761 681 778
rect 657 744 661 761
rect 678 744 681 761
rect 657 727 681 744
rect 657 710 661 727
rect 678 710 681 727
rect 657 693 681 710
rect 657 676 661 693
rect 678 676 681 693
rect 657 659 681 676
rect 657 642 661 659
rect 678 642 681 659
rect 657 625 681 642
rect 657 608 661 625
rect 678 608 681 625
rect 657 591 681 608
rect 657 574 661 591
rect 678 574 681 591
rect 657 557 681 574
rect 657 540 661 557
rect 678 540 681 557
rect 657 523 681 540
rect 657 506 661 523
rect 678 506 681 523
rect 657 489 681 506
rect 657 472 661 489
rect 678 472 681 489
rect 657 455 681 472
rect 657 438 661 455
rect 678 438 681 455
rect 657 421 681 438
rect 657 404 661 421
rect 678 404 681 421
rect 657 387 681 404
rect 657 370 661 387
rect 678 370 681 387
rect 657 353 681 370
rect 657 336 661 353
rect 678 336 681 353
rect 657 319 681 336
rect 657 302 661 319
rect 678 302 681 319
rect 657 285 681 302
rect 657 268 661 285
rect 678 268 681 285
rect 657 251 681 268
rect 657 234 661 251
rect 678 234 681 251
rect 657 217 681 234
rect 657 200 661 217
rect 678 200 681 217
rect 657 183 681 200
rect 657 166 661 183
rect 678 166 681 183
rect 657 158 681 166
rect 702 1137 725 1145
rect 702 1120 705 1137
rect 722 1120 725 1137
rect 702 1103 725 1120
rect 702 1086 705 1103
rect 722 1086 725 1103
rect 702 1069 725 1086
rect 702 1052 705 1069
rect 722 1052 725 1069
rect 702 1035 725 1052
rect 702 1018 705 1035
rect 722 1018 725 1035
rect 702 1001 725 1018
rect 702 984 705 1001
rect 722 984 725 1001
rect 702 967 725 984
rect 702 950 705 967
rect 722 950 725 967
rect 702 933 725 950
rect 702 916 705 933
rect 722 916 725 933
rect 702 899 725 916
rect 702 882 705 899
rect 722 882 725 899
rect 702 865 725 882
rect 702 848 705 865
rect 722 848 725 865
rect 702 831 725 848
rect 702 814 705 831
rect 722 814 725 831
rect 702 797 725 814
rect 702 780 705 797
rect 722 780 725 797
rect 702 763 725 780
rect 702 746 705 763
rect 722 746 725 763
rect 702 729 725 746
rect 702 712 705 729
rect 722 712 725 729
rect 702 695 725 712
rect 702 678 705 695
rect 722 678 725 695
rect 702 661 725 678
rect 702 644 705 661
rect 722 644 725 661
rect 702 627 725 644
rect 702 610 705 627
rect 722 610 725 627
rect 702 593 725 610
rect 702 576 705 593
rect 722 576 725 593
rect 702 559 725 576
rect 702 542 705 559
rect 722 542 725 559
rect 702 525 725 542
rect 702 508 705 525
rect 722 508 725 525
rect 702 491 725 508
rect 702 474 705 491
rect 722 474 725 491
rect 702 457 725 474
rect 702 440 705 457
rect 722 440 725 457
rect 702 423 725 440
rect 702 406 705 423
rect 722 406 725 423
rect 702 389 725 406
rect 702 372 705 389
rect 722 372 725 389
rect 702 355 725 372
rect 702 338 705 355
rect 722 338 725 355
rect 702 321 725 338
rect 702 304 705 321
rect 722 304 725 321
rect 702 287 725 304
rect 702 270 705 287
rect 722 270 725 287
rect 702 253 725 270
rect 702 236 705 253
rect 722 236 725 253
rect 702 219 725 236
rect 702 202 705 219
rect 722 202 725 219
rect 702 185 725 202
rect 702 168 705 185
rect 722 168 725 185
rect 702 115 725 168
rect 746 1135 770 1184
rect 746 1118 749 1135
rect 766 1118 770 1135
rect 746 1101 770 1118
rect 746 1084 749 1101
rect 766 1084 770 1101
rect 746 1067 770 1084
rect 746 1050 749 1067
rect 766 1050 770 1067
rect 746 1033 770 1050
rect 746 1016 749 1033
rect 766 1016 770 1033
rect 746 999 770 1016
rect 746 982 750 999
rect 767 982 770 999
rect 746 965 770 982
rect 746 948 750 965
rect 767 948 770 965
rect 746 931 770 948
rect 746 914 750 931
rect 767 914 770 931
rect 746 897 770 914
rect 746 880 750 897
rect 767 880 770 897
rect 746 863 770 880
rect 746 846 750 863
rect 767 846 770 863
rect 746 829 770 846
rect 746 812 750 829
rect 767 812 770 829
rect 746 795 770 812
rect 746 778 750 795
rect 767 778 770 795
rect 746 761 770 778
rect 746 744 750 761
rect 767 744 770 761
rect 746 727 770 744
rect 746 710 750 727
rect 767 710 770 727
rect 746 693 770 710
rect 746 676 750 693
rect 767 676 770 693
rect 746 659 770 676
rect 746 642 750 659
rect 767 642 770 659
rect 746 625 770 642
rect 746 608 750 625
rect 767 608 770 625
rect 746 591 770 608
rect 746 574 750 591
rect 767 574 770 591
rect 746 557 770 574
rect 746 540 750 557
rect 767 540 770 557
rect 746 523 770 540
rect 746 506 750 523
rect 767 506 770 523
rect 746 489 770 506
rect 746 472 750 489
rect 767 472 770 489
rect 746 455 770 472
rect 746 438 750 455
rect 767 438 770 455
rect 746 421 770 438
rect 746 404 750 421
rect 767 404 770 421
rect 746 387 770 404
rect 746 370 750 387
rect 767 370 770 387
rect 746 353 770 370
rect 746 336 750 353
rect 767 336 770 353
rect 746 319 770 336
rect 746 302 750 319
rect 767 302 770 319
rect 746 285 770 302
rect 746 268 750 285
rect 767 268 770 285
rect 746 251 770 268
rect 746 234 750 251
rect 767 234 770 251
rect 746 217 770 234
rect 746 200 750 217
rect 767 200 770 217
rect 746 183 770 200
rect 746 166 750 183
rect 767 166 770 183
rect 746 158 770 166
rect 791 1135 815 1143
rect 791 1118 794 1135
rect 811 1118 815 1135
rect 791 1101 815 1118
rect 791 1084 794 1101
rect 811 1084 815 1101
rect 791 1067 815 1084
rect 791 1050 794 1067
rect 811 1050 815 1067
rect 791 1033 815 1050
rect 791 1016 794 1033
rect 811 1016 815 1033
rect 791 999 815 1016
rect 791 982 795 999
rect 812 982 815 999
rect 791 965 815 982
rect 791 948 795 965
rect 812 948 815 965
rect 791 931 815 948
rect 791 914 795 931
rect 812 914 815 931
rect 791 897 815 914
rect 791 880 795 897
rect 812 880 815 897
rect 791 863 815 880
rect 791 846 795 863
rect 812 846 815 863
rect 791 829 815 846
rect 791 812 795 829
rect 812 812 815 829
rect 791 795 815 812
rect 791 778 795 795
rect 812 778 815 795
rect 791 761 815 778
rect 791 744 795 761
rect 812 744 815 761
rect 791 727 815 744
rect 791 710 795 727
rect 812 710 815 727
rect 791 693 815 710
rect 791 676 795 693
rect 812 676 815 693
rect 791 659 815 676
rect 791 642 795 659
rect 812 642 815 659
rect 791 625 815 642
rect 791 608 795 625
rect 812 608 815 625
rect 791 591 815 608
rect 791 574 795 591
rect 812 574 815 591
rect 791 557 815 574
rect 791 540 795 557
rect 812 540 815 557
rect 791 523 815 540
rect 791 506 795 523
rect 812 506 815 523
rect 791 489 815 506
rect 791 472 795 489
rect 812 472 815 489
rect 791 455 815 472
rect 791 438 795 455
rect 812 438 815 455
rect 791 421 815 438
rect 791 404 795 421
rect 812 404 815 421
rect 791 387 815 404
rect 791 370 795 387
rect 812 370 815 387
rect 791 353 815 370
rect 791 336 795 353
rect 812 336 815 353
rect 791 319 815 336
rect 791 302 795 319
rect 812 302 815 319
rect 791 285 815 302
rect 791 268 795 285
rect 812 268 815 285
rect 791 251 815 268
rect 791 234 795 251
rect 812 234 815 251
rect 791 217 815 234
rect 791 200 795 217
rect 812 200 815 217
rect 791 183 815 200
rect 791 166 795 183
rect 812 166 815 183
rect 791 115 815 166
rect 836 1135 860 1184
rect 836 1118 839 1135
rect 856 1118 860 1135
rect 836 1101 860 1118
rect 836 1084 839 1101
rect 856 1084 860 1101
rect 836 1067 860 1084
rect 836 1050 839 1067
rect 856 1050 860 1067
rect 836 1033 860 1050
rect 836 1016 839 1033
rect 856 1016 860 1033
rect 836 999 860 1016
rect 836 982 840 999
rect 857 982 860 999
rect 836 965 860 982
rect 836 948 840 965
rect 857 948 860 965
rect 836 931 860 948
rect 836 914 840 931
rect 857 914 860 931
rect 836 897 860 914
rect 836 880 840 897
rect 857 880 860 897
rect 836 863 860 880
rect 836 846 840 863
rect 857 846 860 863
rect 836 829 860 846
rect 836 812 840 829
rect 857 812 860 829
rect 836 795 860 812
rect 836 778 840 795
rect 857 778 860 795
rect 836 761 860 778
rect 836 744 840 761
rect 857 744 860 761
rect 836 727 860 744
rect 836 710 840 727
rect 857 710 860 727
rect 836 693 860 710
rect 836 676 840 693
rect 857 676 860 693
rect 836 659 860 676
rect 836 642 840 659
rect 857 642 860 659
rect 836 625 860 642
rect 836 608 840 625
rect 857 608 860 625
rect 836 591 860 608
rect 836 574 840 591
rect 857 574 860 591
rect 836 557 860 574
rect 836 540 840 557
rect 857 540 860 557
rect 836 523 860 540
rect 836 506 840 523
rect 857 506 860 523
rect 836 489 860 506
rect 836 472 840 489
rect 857 472 860 489
rect 836 455 860 472
rect 836 438 840 455
rect 857 438 860 455
rect 836 421 860 438
rect 836 404 840 421
rect 857 404 860 421
rect 836 387 860 404
rect 836 370 840 387
rect 857 370 860 387
rect 836 353 860 370
rect 836 336 840 353
rect 857 336 860 353
rect 836 319 860 336
rect 836 302 840 319
rect 857 302 860 319
rect 836 285 860 302
rect 836 268 840 285
rect 857 268 860 285
rect 836 251 860 268
rect 836 234 840 251
rect 857 234 860 251
rect 836 217 860 234
rect 836 200 840 217
rect 857 200 860 217
rect 836 183 860 200
rect 836 166 840 183
rect 857 166 860 183
rect 836 158 860 166
rect 881 1135 905 1143
rect 881 1118 884 1135
rect 901 1118 905 1135
rect 881 1101 905 1118
rect 881 1084 884 1101
rect 901 1084 905 1101
rect 881 1067 905 1084
rect 881 1050 884 1067
rect 901 1050 905 1067
rect 881 1033 905 1050
rect 881 1016 884 1033
rect 901 1016 905 1033
rect 881 999 905 1016
rect 881 982 885 999
rect 902 982 905 999
rect 881 965 905 982
rect 881 948 885 965
rect 902 948 905 965
rect 881 931 905 948
rect 881 914 885 931
rect 902 914 905 931
rect 881 897 905 914
rect 881 880 885 897
rect 902 880 905 897
rect 881 863 905 880
rect 881 846 885 863
rect 902 846 905 863
rect 881 829 905 846
rect 881 812 885 829
rect 902 812 905 829
rect 881 795 905 812
rect 881 778 885 795
rect 902 778 905 795
rect 881 761 905 778
rect 881 744 885 761
rect 902 744 905 761
rect 881 727 905 744
rect 881 710 885 727
rect 902 710 905 727
rect 881 693 905 710
rect 881 676 885 693
rect 902 676 905 693
rect 881 659 905 676
rect 881 642 885 659
rect 902 642 905 659
rect 881 625 905 642
rect 881 608 885 625
rect 902 608 905 625
rect 881 591 905 608
rect 881 574 885 591
rect 902 574 905 591
rect 881 557 905 574
rect 881 540 885 557
rect 902 540 905 557
rect 881 523 905 540
rect 881 506 885 523
rect 902 506 905 523
rect 881 489 905 506
rect 881 472 885 489
rect 902 472 905 489
rect 881 455 905 472
rect 881 438 885 455
rect 902 438 905 455
rect 881 421 905 438
rect 881 404 885 421
rect 902 404 905 421
rect 881 387 905 404
rect 881 370 885 387
rect 902 370 905 387
rect 881 353 905 370
rect 881 336 885 353
rect 902 336 905 353
rect 881 319 905 336
rect 881 302 885 319
rect 902 302 905 319
rect 881 285 905 302
rect 881 268 885 285
rect 902 268 905 285
rect 881 251 905 268
rect 881 234 885 251
rect 902 234 905 251
rect 881 217 905 234
rect 881 200 885 217
rect 902 200 905 217
rect 881 183 905 200
rect 881 166 885 183
rect 902 166 905 183
rect 881 115 905 166
rect 926 1135 950 1184
rect 926 1118 929 1135
rect 946 1118 950 1135
rect 926 1101 950 1118
rect 926 1084 929 1101
rect 946 1084 950 1101
rect 926 1067 950 1084
rect 926 1050 929 1067
rect 946 1050 950 1067
rect 926 1033 950 1050
rect 926 1016 929 1033
rect 946 1016 950 1033
rect 926 999 950 1016
rect 926 982 930 999
rect 947 982 950 999
rect 926 965 950 982
rect 926 948 930 965
rect 947 948 950 965
rect 926 931 950 948
rect 926 914 930 931
rect 947 914 950 931
rect 926 897 950 914
rect 926 880 930 897
rect 947 880 950 897
rect 926 863 950 880
rect 926 846 930 863
rect 947 846 950 863
rect 926 829 950 846
rect 926 812 930 829
rect 947 812 950 829
rect 926 795 950 812
rect 926 778 930 795
rect 947 778 950 795
rect 926 761 950 778
rect 926 744 930 761
rect 947 744 950 761
rect 926 727 950 744
rect 926 710 930 727
rect 947 710 950 727
rect 926 693 950 710
rect 926 676 930 693
rect 947 676 950 693
rect 926 659 950 676
rect 926 642 930 659
rect 947 642 950 659
rect 926 625 950 642
rect 926 608 930 625
rect 947 608 950 625
rect 926 591 950 608
rect 926 574 930 591
rect 947 574 950 591
rect 926 557 950 574
rect 926 540 930 557
rect 947 540 950 557
rect 926 523 950 540
rect 926 506 930 523
rect 947 506 950 523
rect 926 489 950 506
rect 926 472 930 489
rect 947 472 950 489
rect 926 455 950 472
rect 926 438 930 455
rect 947 438 950 455
rect 926 421 950 438
rect 926 404 930 421
rect 947 404 950 421
rect 926 387 950 404
rect 926 370 930 387
rect 947 370 950 387
rect 926 353 950 370
rect 926 336 930 353
rect 947 336 950 353
rect 926 319 950 336
rect 926 302 930 319
rect 947 302 950 319
rect 926 285 950 302
rect 926 268 930 285
rect 947 268 950 285
rect 926 251 950 268
rect 926 234 930 251
rect 947 234 950 251
rect 926 217 950 234
rect 926 200 930 217
rect 947 200 950 217
rect 926 183 950 200
rect 926 166 930 183
rect 947 166 950 183
rect 926 158 950 166
rect 971 1135 995 1143
rect 971 1118 974 1135
rect 991 1118 995 1135
rect 971 1101 995 1118
rect 971 1084 974 1101
rect 991 1084 995 1101
rect 971 1067 995 1084
rect 971 1050 974 1067
rect 991 1050 995 1067
rect 971 1033 995 1050
rect 971 1016 974 1033
rect 991 1016 995 1033
rect 971 999 995 1016
rect 971 982 975 999
rect 992 982 995 999
rect 971 965 995 982
rect 971 948 975 965
rect 992 948 995 965
rect 971 931 995 948
rect 971 914 975 931
rect 992 914 995 931
rect 971 897 995 914
rect 971 880 975 897
rect 992 880 995 897
rect 971 863 995 880
rect 971 846 975 863
rect 992 846 995 863
rect 971 829 995 846
rect 971 812 975 829
rect 992 812 995 829
rect 971 795 995 812
rect 971 778 975 795
rect 992 778 995 795
rect 971 761 995 778
rect 971 744 975 761
rect 992 744 995 761
rect 971 727 995 744
rect 971 710 975 727
rect 992 710 995 727
rect 971 693 995 710
rect 971 676 975 693
rect 992 676 995 693
rect 971 659 995 676
rect 971 642 975 659
rect 992 642 995 659
rect 971 625 995 642
rect 971 608 975 625
rect 992 608 995 625
rect 971 591 995 608
rect 971 574 975 591
rect 992 574 995 591
rect 971 557 995 574
rect 971 540 975 557
rect 992 540 995 557
rect 971 523 995 540
rect 971 506 975 523
rect 992 506 995 523
rect 971 489 995 506
rect 971 472 975 489
rect 992 472 995 489
rect 971 455 995 472
rect 971 438 975 455
rect 992 438 995 455
rect 971 421 995 438
rect 971 404 975 421
rect 992 404 995 421
rect 971 387 995 404
rect 971 370 975 387
rect 992 370 995 387
rect 971 353 995 370
rect 971 336 975 353
rect 992 336 995 353
rect 971 319 995 336
rect 971 302 975 319
rect 992 302 995 319
rect 971 285 995 302
rect 971 268 975 285
rect 992 268 995 285
rect 971 251 995 268
rect 971 234 975 251
rect 992 234 995 251
rect 971 217 995 234
rect 971 200 975 217
rect 992 200 995 217
rect 971 183 995 200
rect 971 166 975 183
rect 992 166 995 183
rect 971 115 995 166
rect 1017 1135 1041 1184
rect 1017 1118 1020 1135
rect 1037 1118 1041 1135
rect 1017 1101 1041 1118
rect 1017 1084 1020 1101
rect 1037 1084 1041 1101
rect 1017 1067 1041 1084
rect 1017 1050 1020 1067
rect 1037 1050 1041 1067
rect 1017 1033 1041 1050
rect 1017 1016 1020 1033
rect 1037 1016 1041 1033
rect 1017 999 1041 1016
rect 1017 982 1021 999
rect 1038 982 1041 999
rect 1017 965 1041 982
rect 1017 948 1021 965
rect 1038 948 1041 965
rect 1017 931 1041 948
rect 1017 914 1021 931
rect 1038 914 1041 931
rect 1017 897 1041 914
rect 1017 880 1021 897
rect 1038 880 1041 897
rect 1017 863 1041 880
rect 1017 846 1021 863
rect 1038 846 1041 863
rect 1017 829 1041 846
rect 1017 812 1021 829
rect 1038 812 1041 829
rect 1017 795 1041 812
rect 1017 778 1021 795
rect 1038 778 1041 795
rect 1017 761 1041 778
rect 1017 744 1021 761
rect 1038 744 1041 761
rect 1017 727 1041 744
rect 1017 710 1021 727
rect 1038 710 1041 727
rect 1017 693 1041 710
rect 1017 676 1021 693
rect 1038 676 1041 693
rect 1017 659 1041 676
rect 1017 642 1021 659
rect 1038 642 1041 659
rect 1017 625 1041 642
rect 1017 608 1021 625
rect 1038 608 1041 625
rect 1017 591 1041 608
rect 1017 574 1021 591
rect 1038 574 1041 591
rect 1017 557 1041 574
rect 1017 540 1021 557
rect 1038 540 1041 557
rect 1017 523 1041 540
rect 1017 506 1021 523
rect 1038 506 1041 523
rect 1017 489 1041 506
rect 1017 472 1021 489
rect 1038 472 1041 489
rect 1017 455 1041 472
rect 1017 438 1021 455
rect 1038 438 1041 455
rect 1017 421 1041 438
rect 1017 404 1021 421
rect 1038 404 1041 421
rect 1017 387 1041 404
rect 1017 370 1021 387
rect 1038 370 1041 387
rect 1017 353 1041 370
rect 1017 336 1021 353
rect 1038 336 1041 353
rect 1017 319 1041 336
rect 1017 302 1021 319
rect 1038 302 1041 319
rect 1017 285 1041 302
rect 1017 268 1021 285
rect 1038 268 1041 285
rect 1017 251 1041 268
rect 1017 234 1021 251
rect 1038 234 1041 251
rect 1017 217 1041 234
rect 1017 200 1021 217
rect 1038 200 1041 217
rect 1017 183 1041 200
rect 1017 166 1021 183
rect 1038 166 1041 183
rect 1017 158 1041 166
rect 1062 1137 1085 1145
rect 1062 1120 1065 1137
rect 1082 1120 1085 1137
rect 1062 1103 1085 1120
rect 1062 1086 1065 1103
rect 1082 1086 1085 1103
rect 1062 1069 1085 1086
rect 1062 1052 1065 1069
rect 1082 1052 1085 1069
rect 1062 1035 1085 1052
rect 1062 1018 1065 1035
rect 1082 1018 1085 1035
rect 1062 1001 1085 1018
rect 1062 984 1065 1001
rect 1082 984 1085 1001
rect 1062 967 1085 984
rect 1062 950 1065 967
rect 1082 950 1085 967
rect 1062 933 1085 950
rect 1062 916 1065 933
rect 1082 916 1085 933
rect 1062 899 1085 916
rect 1062 882 1065 899
rect 1082 882 1085 899
rect 1062 865 1085 882
rect 1062 848 1065 865
rect 1082 848 1085 865
rect 1062 831 1085 848
rect 1062 814 1065 831
rect 1082 814 1085 831
rect 1062 797 1085 814
rect 1062 780 1065 797
rect 1082 780 1085 797
rect 1062 763 1085 780
rect 1062 746 1065 763
rect 1082 746 1085 763
rect 1062 729 1085 746
rect 1062 712 1065 729
rect 1082 712 1085 729
rect 1062 695 1085 712
rect 1062 678 1065 695
rect 1082 678 1085 695
rect 1062 661 1085 678
rect 1062 644 1065 661
rect 1082 644 1085 661
rect 1062 627 1085 644
rect 1062 610 1065 627
rect 1082 610 1085 627
rect 1062 593 1085 610
rect 1062 576 1065 593
rect 1082 576 1085 593
rect 1062 559 1085 576
rect 1062 542 1065 559
rect 1082 542 1085 559
rect 1062 525 1085 542
rect 1062 508 1065 525
rect 1082 508 1085 525
rect 1062 491 1085 508
rect 1062 474 1065 491
rect 1082 474 1085 491
rect 1062 457 1085 474
rect 1062 440 1065 457
rect 1082 440 1085 457
rect 1062 423 1085 440
rect 1062 406 1065 423
rect 1082 406 1085 423
rect 1062 389 1085 406
rect 1062 372 1065 389
rect 1082 372 1085 389
rect 1062 355 1085 372
rect 1062 338 1065 355
rect 1082 338 1085 355
rect 1062 321 1085 338
rect 1062 304 1065 321
rect 1082 304 1085 321
rect 1062 287 1085 304
rect 1062 270 1065 287
rect 1082 270 1085 287
rect 1062 253 1085 270
rect 1062 236 1065 253
rect 1082 236 1085 253
rect 1062 219 1085 236
rect 1062 202 1065 219
rect 1082 202 1085 219
rect 1062 185 1085 202
rect 1062 168 1065 185
rect 1082 168 1085 185
rect 1062 115 1085 168
rect 1106 1135 1130 1184
rect 1106 1118 1109 1135
rect 1126 1118 1130 1135
rect 1106 1101 1130 1118
rect 1106 1084 1109 1101
rect 1126 1084 1130 1101
rect 1106 1067 1130 1084
rect 1106 1050 1109 1067
rect 1126 1050 1130 1067
rect 1106 1033 1130 1050
rect 1106 1016 1109 1033
rect 1126 1016 1130 1033
rect 1106 999 1130 1016
rect 1106 982 1110 999
rect 1127 982 1130 999
rect 1106 965 1130 982
rect 1106 948 1110 965
rect 1127 948 1130 965
rect 1106 931 1130 948
rect 1106 914 1110 931
rect 1127 914 1130 931
rect 1106 897 1130 914
rect 1106 880 1110 897
rect 1127 880 1130 897
rect 1106 863 1130 880
rect 1106 846 1110 863
rect 1127 846 1130 863
rect 1106 829 1130 846
rect 1106 812 1110 829
rect 1127 812 1130 829
rect 1106 795 1130 812
rect 1106 778 1110 795
rect 1127 778 1130 795
rect 1106 761 1130 778
rect 1106 744 1110 761
rect 1127 744 1130 761
rect 1106 727 1130 744
rect 1106 710 1110 727
rect 1127 710 1130 727
rect 1106 693 1130 710
rect 1106 676 1110 693
rect 1127 676 1130 693
rect 1106 659 1130 676
rect 1106 642 1110 659
rect 1127 642 1130 659
rect 1106 625 1130 642
rect 1106 608 1110 625
rect 1127 608 1130 625
rect 1106 591 1130 608
rect 1106 574 1110 591
rect 1127 574 1130 591
rect 1106 557 1130 574
rect 1106 540 1110 557
rect 1127 540 1130 557
rect 1106 523 1130 540
rect 1106 506 1110 523
rect 1127 506 1130 523
rect 1106 489 1130 506
rect 1106 472 1110 489
rect 1127 472 1130 489
rect 1106 455 1130 472
rect 1106 438 1110 455
rect 1127 438 1130 455
rect 1106 421 1130 438
rect 1106 404 1110 421
rect 1127 404 1130 421
rect 1106 387 1130 404
rect 1106 370 1110 387
rect 1127 370 1130 387
rect 1106 353 1130 370
rect 1106 336 1110 353
rect 1127 336 1130 353
rect 1106 319 1130 336
rect 1106 302 1110 319
rect 1127 302 1130 319
rect 1106 285 1130 302
rect 1106 268 1110 285
rect 1127 268 1130 285
rect 1106 251 1130 268
rect 1106 234 1110 251
rect 1127 234 1130 251
rect 1106 217 1130 234
rect 1106 200 1110 217
rect 1127 200 1130 217
rect 1106 183 1130 200
rect 1106 166 1110 183
rect 1127 166 1130 183
rect 1106 158 1130 166
rect 1151 1135 1175 1143
rect 1151 1118 1154 1135
rect 1171 1118 1175 1135
rect 1151 1101 1175 1118
rect 1151 1084 1154 1101
rect 1171 1084 1175 1101
rect 1151 1067 1175 1084
rect 1151 1050 1154 1067
rect 1171 1050 1175 1067
rect 1151 1033 1175 1050
rect 1151 1016 1154 1033
rect 1171 1016 1175 1033
rect 1151 999 1175 1016
rect 1151 982 1155 999
rect 1172 982 1175 999
rect 1151 965 1175 982
rect 1151 948 1155 965
rect 1172 948 1175 965
rect 1151 931 1175 948
rect 1151 914 1155 931
rect 1172 914 1175 931
rect 1151 897 1175 914
rect 1151 880 1155 897
rect 1172 880 1175 897
rect 1151 863 1175 880
rect 1151 846 1155 863
rect 1172 846 1175 863
rect 1151 829 1175 846
rect 1151 812 1155 829
rect 1172 812 1175 829
rect 1151 795 1175 812
rect 1151 778 1155 795
rect 1172 778 1175 795
rect 1151 761 1175 778
rect 1151 744 1155 761
rect 1172 744 1175 761
rect 1151 727 1175 744
rect 1151 710 1155 727
rect 1172 710 1175 727
rect 1151 693 1175 710
rect 1151 676 1155 693
rect 1172 676 1175 693
rect 1151 659 1175 676
rect 1151 642 1155 659
rect 1172 642 1175 659
rect 1151 625 1175 642
rect 1151 608 1155 625
rect 1172 608 1175 625
rect 1151 591 1175 608
rect 1151 574 1155 591
rect 1172 574 1175 591
rect 1151 557 1175 574
rect 1151 540 1155 557
rect 1172 540 1175 557
rect 1151 523 1175 540
rect 1151 506 1155 523
rect 1172 506 1175 523
rect 1151 489 1175 506
rect 1151 472 1155 489
rect 1172 472 1175 489
rect 1151 455 1175 472
rect 1151 438 1155 455
rect 1172 438 1175 455
rect 1151 421 1175 438
rect 1151 404 1155 421
rect 1172 404 1175 421
rect 1151 387 1175 404
rect 1151 370 1155 387
rect 1172 370 1175 387
rect 1151 353 1175 370
rect 1151 336 1155 353
rect 1172 336 1175 353
rect 1151 319 1175 336
rect 1151 302 1155 319
rect 1172 302 1175 319
rect 1151 285 1175 302
rect 1151 268 1155 285
rect 1172 268 1175 285
rect 1151 251 1175 268
rect 1151 234 1155 251
rect 1172 234 1175 251
rect 1151 217 1175 234
rect 1151 200 1155 217
rect 1172 200 1175 217
rect 1151 183 1175 200
rect 1151 166 1155 183
rect 1172 166 1175 183
rect 1151 115 1175 166
rect 1196 1135 1220 1184
rect 1196 1118 1199 1135
rect 1216 1118 1220 1135
rect 1196 1101 1220 1118
rect 1196 1084 1199 1101
rect 1216 1084 1220 1101
rect 1196 1067 1220 1084
rect 1196 1050 1199 1067
rect 1216 1050 1220 1067
rect 1196 1033 1220 1050
rect 1196 1016 1199 1033
rect 1216 1016 1220 1033
rect 1196 999 1220 1016
rect 1196 982 1200 999
rect 1217 982 1220 999
rect 1196 965 1220 982
rect 1196 948 1200 965
rect 1217 948 1220 965
rect 1196 931 1220 948
rect 1196 914 1200 931
rect 1217 914 1220 931
rect 1196 897 1220 914
rect 1196 880 1200 897
rect 1217 880 1220 897
rect 1196 863 1220 880
rect 1196 846 1200 863
rect 1217 846 1220 863
rect 1196 829 1220 846
rect 1196 812 1200 829
rect 1217 812 1220 829
rect 1196 795 1220 812
rect 1196 778 1200 795
rect 1217 778 1220 795
rect 1196 761 1220 778
rect 1196 744 1200 761
rect 1217 744 1220 761
rect 1196 727 1220 744
rect 1196 710 1200 727
rect 1217 710 1220 727
rect 1196 693 1220 710
rect 1196 676 1200 693
rect 1217 676 1220 693
rect 1196 659 1220 676
rect 1196 642 1200 659
rect 1217 642 1220 659
rect 1196 625 1220 642
rect 1196 608 1200 625
rect 1217 608 1220 625
rect 1196 591 1220 608
rect 1196 574 1200 591
rect 1217 574 1220 591
rect 1196 557 1220 574
rect 1196 540 1200 557
rect 1217 540 1220 557
rect 1196 523 1220 540
rect 1196 506 1200 523
rect 1217 506 1220 523
rect 1196 489 1220 506
rect 1196 472 1200 489
rect 1217 472 1220 489
rect 1196 455 1220 472
rect 1196 438 1200 455
rect 1217 438 1220 455
rect 1196 421 1220 438
rect 1196 404 1200 421
rect 1217 404 1220 421
rect 1196 387 1220 404
rect 1196 370 1200 387
rect 1217 370 1220 387
rect 1196 353 1220 370
rect 1196 336 1200 353
rect 1217 336 1220 353
rect 1196 319 1220 336
rect 1196 302 1200 319
rect 1217 302 1220 319
rect 1196 285 1220 302
rect 1196 268 1200 285
rect 1217 268 1220 285
rect 1196 251 1220 268
rect 1196 234 1200 251
rect 1217 234 1220 251
rect 1196 217 1220 234
rect 1196 200 1200 217
rect 1217 200 1220 217
rect 1196 183 1220 200
rect 1196 166 1200 183
rect 1217 166 1220 183
rect 1196 158 1220 166
rect 1241 1135 1265 1143
rect 1241 1118 1244 1135
rect 1261 1118 1265 1135
rect 1241 1101 1265 1118
rect 1241 1084 1244 1101
rect 1261 1084 1265 1101
rect 1241 1067 1265 1084
rect 1241 1050 1244 1067
rect 1261 1050 1265 1067
rect 1241 1033 1265 1050
rect 1241 1016 1244 1033
rect 1261 1016 1265 1033
rect 1241 999 1265 1016
rect 1241 982 1245 999
rect 1262 982 1265 999
rect 1241 965 1265 982
rect 1241 948 1245 965
rect 1262 948 1265 965
rect 1241 931 1265 948
rect 1241 914 1245 931
rect 1262 914 1265 931
rect 1241 897 1265 914
rect 1241 880 1245 897
rect 1262 880 1265 897
rect 1241 863 1265 880
rect 1241 846 1245 863
rect 1262 846 1265 863
rect 1241 829 1265 846
rect 1241 812 1245 829
rect 1262 812 1265 829
rect 1241 795 1265 812
rect 1241 778 1245 795
rect 1262 778 1265 795
rect 1241 761 1265 778
rect 1241 744 1245 761
rect 1262 744 1265 761
rect 1241 727 1265 744
rect 1241 710 1245 727
rect 1262 710 1265 727
rect 1241 693 1265 710
rect 1241 676 1245 693
rect 1262 676 1265 693
rect 1241 659 1265 676
rect 1241 642 1245 659
rect 1262 642 1265 659
rect 1241 625 1265 642
rect 1241 608 1245 625
rect 1262 608 1265 625
rect 1241 591 1265 608
rect 1241 574 1245 591
rect 1262 574 1265 591
rect 1241 557 1265 574
rect 1241 540 1245 557
rect 1262 540 1265 557
rect 1241 523 1265 540
rect 1241 506 1245 523
rect 1262 506 1265 523
rect 1241 489 1265 506
rect 1241 472 1245 489
rect 1262 472 1265 489
rect 1241 455 1265 472
rect 1241 438 1245 455
rect 1262 438 1265 455
rect 1241 421 1265 438
rect 1241 404 1245 421
rect 1262 404 1265 421
rect 1241 387 1265 404
rect 1241 370 1245 387
rect 1262 370 1265 387
rect 1241 353 1265 370
rect 1241 336 1245 353
rect 1262 336 1265 353
rect 1241 319 1265 336
rect 1241 302 1245 319
rect 1262 302 1265 319
rect 1241 285 1265 302
rect 1241 268 1245 285
rect 1262 268 1265 285
rect 1241 251 1265 268
rect 1241 234 1245 251
rect 1262 234 1265 251
rect 1241 217 1265 234
rect 1241 200 1245 217
rect 1262 200 1265 217
rect 1241 183 1265 200
rect 1241 166 1245 183
rect 1262 166 1265 183
rect 1241 115 1265 166
rect 1286 1135 1310 1184
rect 1286 1118 1289 1135
rect 1306 1118 1310 1135
rect 1286 1101 1310 1118
rect 1286 1084 1289 1101
rect 1306 1084 1310 1101
rect 1286 1067 1310 1084
rect 1286 1050 1289 1067
rect 1306 1050 1310 1067
rect 1286 1033 1310 1050
rect 1286 1016 1289 1033
rect 1306 1016 1310 1033
rect 1286 999 1310 1016
rect 1286 982 1290 999
rect 1307 982 1310 999
rect 1286 965 1310 982
rect 1286 948 1290 965
rect 1307 948 1310 965
rect 1286 931 1310 948
rect 1286 914 1290 931
rect 1307 914 1310 931
rect 1286 897 1310 914
rect 1286 880 1290 897
rect 1307 880 1310 897
rect 1286 863 1310 880
rect 1286 846 1290 863
rect 1307 846 1310 863
rect 1286 829 1310 846
rect 1286 812 1290 829
rect 1307 812 1310 829
rect 1286 795 1310 812
rect 1286 778 1290 795
rect 1307 778 1310 795
rect 1286 761 1310 778
rect 1286 744 1290 761
rect 1307 744 1310 761
rect 1286 727 1310 744
rect 1286 710 1290 727
rect 1307 710 1310 727
rect 1286 693 1310 710
rect 1286 676 1290 693
rect 1307 676 1310 693
rect 1286 659 1310 676
rect 1286 642 1290 659
rect 1307 642 1310 659
rect 1286 625 1310 642
rect 1286 608 1290 625
rect 1307 608 1310 625
rect 1286 591 1310 608
rect 1286 574 1290 591
rect 1307 574 1310 591
rect 1286 557 1310 574
rect 1286 540 1290 557
rect 1307 540 1310 557
rect 1286 523 1310 540
rect 1286 506 1290 523
rect 1307 506 1310 523
rect 1286 489 1310 506
rect 1286 472 1290 489
rect 1307 472 1310 489
rect 1286 455 1310 472
rect 1286 438 1290 455
rect 1307 438 1310 455
rect 1286 421 1310 438
rect 1286 404 1290 421
rect 1307 404 1310 421
rect 1286 387 1310 404
rect 1286 370 1290 387
rect 1307 370 1310 387
rect 1286 353 1310 370
rect 1286 336 1290 353
rect 1307 336 1310 353
rect 1286 319 1310 336
rect 1286 302 1290 319
rect 1307 302 1310 319
rect 1286 285 1310 302
rect 1286 268 1290 285
rect 1307 268 1310 285
rect 1286 251 1310 268
rect 1286 234 1290 251
rect 1307 234 1310 251
rect 1286 217 1310 234
rect 1286 200 1290 217
rect 1307 200 1310 217
rect 1286 183 1310 200
rect 1286 166 1290 183
rect 1307 166 1310 183
rect 1286 158 1310 166
rect 1331 1135 1355 1143
rect 1331 1118 1334 1135
rect 1351 1118 1355 1135
rect 1331 1101 1355 1118
rect 1331 1084 1334 1101
rect 1351 1084 1355 1101
rect 1331 1067 1355 1084
rect 1331 1050 1334 1067
rect 1351 1050 1355 1067
rect 1331 1033 1355 1050
rect 1331 1016 1334 1033
rect 1351 1016 1355 1033
rect 1331 999 1355 1016
rect 1331 982 1335 999
rect 1352 982 1355 999
rect 1331 965 1355 982
rect 1331 948 1335 965
rect 1352 948 1355 965
rect 1331 931 1355 948
rect 1331 914 1335 931
rect 1352 914 1355 931
rect 1331 897 1355 914
rect 1331 880 1335 897
rect 1352 880 1355 897
rect 1331 863 1355 880
rect 1331 846 1335 863
rect 1352 846 1355 863
rect 1331 829 1355 846
rect 1331 812 1335 829
rect 1352 812 1355 829
rect 1331 795 1355 812
rect 1331 778 1335 795
rect 1352 778 1355 795
rect 1331 761 1355 778
rect 1331 744 1335 761
rect 1352 744 1355 761
rect 1331 727 1355 744
rect 1331 710 1335 727
rect 1352 710 1355 727
rect 1331 693 1355 710
rect 1331 676 1335 693
rect 1352 676 1355 693
rect 1331 659 1355 676
rect 1331 642 1335 659
rect 1352 642 1355 659
rect 1331 625 1355 642
rect 1331 608 1335 625
rect 1352 608 1355 625
rect 1331 591 1355 608
rect 1331 574 1335 591
rect 1352 574 1355 591
rect 1331 557 1355 574
rect 1331 540 1335 557
rect 1352 540 1355 557
rect 1331 523 1355 540
rect 1331 506 1335 523
rect 1352 506 1355 523
rect 1331 489 1355 506
rect 1331 472 1335 489
rect 1352 472 1355 489
rect 1331 455 1355 472
rect 1331 438 1335 455
rect 1352 438 1355 455
rect 1331 421 1355 438
rect 1331 404 1335 421
rect 1352 404 1355 421
rect 1331 387 1355 404
rect 1331 370 1335 387
rect 1352 370 1355 387
rect 1331 353 1355 370
rect 1331 336 1335 353
rect 1352 336 1355 353
rect 1331 319 1355 336
rect 1331 302 1335 319
rect 1352 302 1355 319
rect 1331 285 1355 302
rect 1331 268 1335 285
rect 1352 268 1355 285
rect 1331 251 1355 268
rect 1331 234 1335 251
rect 1352 234 1355 251
rect 1331 217 1355 234
rect 1331 200 1335 217
rect 1352 200 1355 217
rect 1331 183 1355 200
rect 1331 166 1335 183
rect 1352 166 1355 183
rect 1331 115 1355 166
rect 1376 1135 1400 1184
rect 1376 1118 1379 1135
rect 1396 1118 1400 1135
rect 1376 1101 1400 1118
rect 1376 1084 1379 1101
rect 1396 1084 1400 1101
rect 1376 1067 1400 1084
rect 1376 1050 1379 1067
rect 1396 1050 1400 1067
rect 1376 1033 1400 1050
rect 1376 1016 1379 1033
rect 1396 1016 1400 1033
rect 1376 999 1400 1016
rect 1376 982 1380 999
rect 1397 982 1400 999
rect 1376 965 1400 982
rect 1376 948 1380 965
rect 1397 948 1400 965
rect 1376 931 1400 948
rect 1376 914 1380 931
rect 1397 914 1400 931
rect 1376 897 1400 914
rect 1376 880 1380 897
rect 1397 880 1400 897
rect 1376 863 1400 880
rect 1376 846 1380 863
rect 1397 846 1400 863
rect 1376 829 1400 846
rect 1376 812 1380 829
rect 1397 812 1400 829
rect 1376 795 1400 812
rect 1376 778 1380 795
rect 1397 778 1400 795
rect 1376 761 1400 778
rect 1376 744 1380 761
rect 1397 744 1400 761
rect 1376 727 1400 744
rect 1376 710 1380 727
rect 1397 710 1400 727
rect 1376 693 1400 710
rect 1376 676 1380 693
rect 1397 676 1400 693
rect 1376 659 1400 676
rect 1376 642 1380 659
rect 1397 642 1400 659
rect 1376 625 1400 642
rect 1376 608 1380 625
rect 1397 608 1400 625
rect 1376 591 1400 608
rect 1376 574 1380 591
rect 1397 574 1400 591
rect 1376 557 1400 574
rect 1376 540 1380 557
rect 1397 540 1400 557
rect 1376 523 1400 540
rect 1376 506 1380 523
rect 1397 506 1400 523
rect 1376 489 1400 506
rect 1376 472 1380 489
rect 1397 472 1400 489
rect 1376 455 1400 472
rect 1376 438 1380 455
rect 1397 438 1400 455
rect 1376 421 1400 438
rect 1376 404 1380 421
rect 1397 404 1400 421
rect 1376 387 1400 404
rect 1376 370 1380 387
rect 1397 370 1400 387
rect 1376 353 1400 370
rect 1376 336 1380 353
rect 1397 336 1400 353
rect 1376 319 1400 336
rect 1376 302 1380 319
rect 1397 302 1400 319
rect 1376 285 1400 302
rect 1376 268 1380 285
rect 1397 268 1400 285
rect 1376 251 1400 268
rect 1376 234 1380 251
rect 1397 234 1400 251
rect 1376 217 1400 234
rect 1376 200 1380 217
rect 1397 200 1400 217
rect 1376 183 1400 200
rect 1376 166 1380 183
rect 1397 166 1400 183
rect 1376 158 1400 166
rect 1421 1137 1444 1145
rect 1421 1120 1424 1137
rect 1441 1120 1444 1137
rect 1421 1103 1444 1120
rect 1421 1086 1424 1103
rect 1441 1086 1444 1103
rect 1421 1069 1444 1086
rect 1421 1052 1424 1069
rect 1441 1052 1444 1069
rect 1421 1035 1444 1052
rect 1421 1018 1424 1035
rect 1441 1018 1444 1035
rect 1421 1001 1444 1018
rect 1421 984 1424 1001
rect 1441 984 1444 1001
rect 1421 967 1444 984
rect 1421 950 1424 967
rect 1441 950 1444 967
rect 1421 933 1444 950
rect 1421 916 1424 933
rect 1441 916 1444 933
rect 1421 899 1444 916
rect 1421 882 1424 899
rect 1441 882 1444 899
rect 1421 865 1444 882
rect 1421 848 1424 865
rect 1441 848 1444 865
rect 1421 831 1444 848
rect 1421 814 1424 831
rect 1441 814 1444 831
rect 1421 797 1444 814
rect 1421 780 1424 797
rect 1441 780 1444 797
rect 1421 763 1444 780
rect 1421 746 1424 763
rect 1441 746 1444 763
rect 1421 729 1444 746
rect 1421 712 1424 729
rect 1441 712 1444 729
rect 1421 695 1444 712
rect 1421 678 1424 695
rect 1441 678 1444 695
rect 1421 661 1444 678
rect 1421 644 1424 661
rect 1441 644 1444 661
rect 1421 627 1444 644
rect 1421 610 1424 627
rect 1441 610 1444 627
rect 1421 593 1444 610
rect 1421 576 1424 593
rect 1441 576 1444 593
rect 1421 559 1444 576
rect 1421 542 1424 559
rect 1441 542 1444 559
rect 1421 525 1444 542
rect 1421 508 1424 525
rect 1441 508 1444 525
rect 1421 491 1444 508
rect 1421 474 1424 491
rect 1441 474 1444 491
rect 1421 457 1444 474
rect 1421 440 1424 457
rect 1441 440 1444 457
rect 1421 423 1444 440
rect 1421 406 1424 423
rect 1441 406 1444 423
rect 1421 389 1444 406
rect 1421 372 1424 389
rect 1441 372 1444 389
rect 1421 355 1444 372
rect 1421 338 1424 355
rect 1441 338 1444 355
rect 1421 321 1444 338
rect 1421 304 1424 321
rect 1441 304 1444 321
rect 1421 287 1444 304
rect 1421 270 1424 287
rect 1441 270 1444 287
rect 1421 253 1444 270
rect 1421 236 1424 253
rect 1441 236 1444 253
rect 1421 219 1444 236
rect 1421 202 1424 219
rect 1441 202 1444 219
rect 1421 185 1444 202
rect 1421 168 1424 185
rect 1441 168 1444 185
rect 1421 115 1444 168
rect 1465 1135 1489 1184
rect 1465 1118 1468 1135
rect 1485 1118 1489 1135
rect 1465 1101 1489 1118
rect 1465 1084 1468 1101
rect 1485 1084 1489 1101
rect 1465 1067 1489 1084
rect 1465 1050 1468 1067
rect 1485 1050 1489 1067
rect 1465 1033 1489 1050
rect 1465 1016 1468 1033
rect 1485 1016 1489 1033
rect 1465 999 1489 1016
rect 1465 982 1469 999
rect 1486 982 1489 999
rect 1465 965 1489 982
rect 1465 948 1469 965
rect 1486 948 1489 965
rect 1465 931 1489 948
rect 1465 914 1469 931
rect 1486 914 1489 931
rect 1465 897 1489 914
rect 1465 880 1469 897
rect 1486 880 1489 897
rect 1465 863 1489 880
rect 1465 846 1469 863
rect 1486 846 1489 863
rect 1465 829 1489 846
rect 1465 812 1469 829
rect 1486 812 1489 829
rect 1465 795 1489 812
rect 1465 778 1469 795
rect 1486 778 1489 795
rect 1465 761 1489 778
rect 1465 744 1469 761
rect 1486 744 1489 761
rect 1465 727 1489 744
rect 1465 710 1469 727
rect 1486 710 1489 727
rect 1465 693 1489 710
rect 1465 676 1469 693
rect 1486 676 1489 693
rect 1465 659 1489 676
rect 1465 642 1469 659
rect 1486 642 1489 659
rect 1465 625 1489 642
rect 1465 608 1469 625
rect 1486 608 1489 625
rect 1465 591 1489 608
rect 1465 574 1469 591
rect 1486 574 1489 591
rect 1465 557 1489 574
rect 1465 540 1469 557
rect 1486 540 1489 557
rect 1465 523 1489 540
rect 1465 506 1469 523
rect 1486 506 1489 523
rect 1465 489 1489 506
rect 1465 472 1469 489
rect 1486 472 1489 489
rect 1465 455 1489 472
rect 1465 438 1469 455
rect 1486 438 1489 455
rect 1465 421 1489 438
rect 1465 404 1469 421
rect 1486 404 1489 421
rect 1465 387 1489 404
rect 1465 370 1469 387
rect 1486 370 1489 387
rect 1465 353 1489 370
rect 1465 336 1469 353
rect 1486 336 1489 353
rect 1465 319 1489 336
rect 1465 302 1469 319
rect 1486 302 1489 319
rect 1465 285 1489 302
rect 1465 268 1469 285
rect 1486 268 1489 285
rect 1465 251 1489 268
rect 1465 234 1469 251
rect 1486 234 1489 251
rect 1465 217 1489 234
rect 1465 200 1469 217
rect 1486 200 1489 217
rect 1465 183 1489 200
rect 1465 166 1469 183
rect 1486 166 1489 183
rect 1465 158 1489 166
rect 1510 1135 1534 1143
rect 1510 1118 1513 1135
rect 1530 1118 1534 1135
rect 1510 1101 1534 1118
rect 1510 1084 1513 1101
rect 1530 1084 1534 1101
rect 1510 1067 1534 1084
rect 1510 1050 1513 1067
rect 1530 1050 1534 1067
rect 1510 1033 1534 1050
rect 1510 1016 1513 1033
rect 1530 1016 1534 1033
rect 1510 999 1534 1016
rect 1510 982 1514 999
rect 1531 982 1534 999
rect 1510 965 1534 982
rect 1510 948 1514 965
rect 1531 948 1534 965
rect 1510 931 1534 948
rect 1510 914 1514 931
rect 1531 914 1534 931
rect 1510 897 1534 914
rect 1510 880 1514 897
rect 1531 880 1534 897
rect 1510 863 1534 880
rect 1510 846 1514 863
rect 1531 846 1534 863
rect 1510 829 1534 846
rect 1510 812 1514 829
rect 1531 812 1534 829
rect 1510 795 1534 812
rect 1510 778 1514 795
rect 1531 778 1534 795
rect 1510 761 1534 778
rect 1510 744 1514 761
rect 1531 744 1534 761
rect 1510 727 1534 744
rect 1510 710 1514 727
rect 1531 710 1534 727
rect 1510 693 1534 710
rect 1510 676 1514 693
rect 1531 676 1534 693
rect 1510 659 1534 676
rect 1510 642 1514 659
rect 1531 642 1534 659
rect 1510 625 1534 642
rect 1510 608 1514 625
rect 1531 608 1534 625
rect 1510 591 1534 608
rect 1510 574 1514 591
rect 1531 574 1534 591
rect 1510 557 1534 574
rect 1510 540 1514 557
rect 1531 540 1534 557
rect 1510 523 1534 540
rect 1510 506 1514 523
rect 1531 506 1534 523
rect 1510 489 1534 506
rect 1510 472 1514 489
rect 1531 472 1534 489
rect 1510 455 1534 472
rect 1510 438 1514 455
rect 1531 438 1534 455
rect 1510 421 1534 438
rect 1510 404 1514 421
rect 1531 404 1534 421
rect 1510 387 1534 404
rect 1510 370 1514 387
rect 1531 370 1534 387
rect 1510 353 1534 370
rect 1510 336 1514 353
rect 1531 336 1534 353
rect 1510 319 1534 336
rect 1510 302 1514 319
rect 1531 302 1534 319
rect 1510 285 1534 302
rect 1510 268 1514 285
rect 1531 268 1534 285
rect 1510 251 1534 268
rect 1510 234 1514 251
rect 1531 234 1534 251
rect 1510 217 1534 234
rect 1510 200 1514 217
rect 1531 200 1534 217
rect 1510 183 1534 200
rect 1510 166 1514 183
rect 1531 166 1534 183
rect 1510 115 1534 166
rect 1555 1135 1579 1184
rect 1555 1118 1558 1135
rect 1575 1118 1579 1135
rect 1555 1101 1579 1118
rect 1555 1084 1558 1101
rect 1575 1084 1579 1101
rect 1555 1067 1579 1084
rect 1555 1050 1558 1067
rect 1575 1050 1579 1067
rect 1555 1033 1579 1050
rect 1555 1016 1558 1033
rect 1575 1016 1579 1033
rect 1555 999 1579 1016
rect 1555 982 1559 999
rect 1576 982 1579 999
rect 1555 965 1579 982
rect 1555 948 1559 965
rect 1576 948 1579 965
rect 1555 931 1579 948
rect 1555 914 1559 931
rect 1576 914 1579 931
rect 1555 897 1579 914
rect 1555 880 1559 897
rect 1576 880 1579 897
rect 1555 863 1579 880
rect 1555 846 1559 863
rect 1576 846 1579 863
rect 1555 829 1579 846
rect 1555 812 1559 829
rect 1576 812 1579 829
rect 1555 795 1579 812
rect 1555 778 1559 795
rect 1576 778 1579 795
rect 1555 761 1579 778
rect 1555 744 1559 761
rect 1576 744 1579 761
rect 1555 727 1579 744
rect 1555 710 1559 727
rect 1576 710 1579 727
rect 1555 693 1579 710
rect 1555 676 1559 693
rect 1576 676 1579 693
rect 1555 659 1579 676
rect 1555 642 1559 659
rect 1576 642 1579 659
rect 1555 625 1579 642
rect 1555 608 1559 625
rect 1576 608 1579 625
rect 1555 591 1579 608
rect 1555 574 1559 591
rect 1576 574 1579 591
rect 1555 557 1579 574
rect 1555 540 1559 557
rect 1576 540 1579 557
rect 1555 523 1579 540
rect 1555 506 1559 523
rect 1576 506 1579 523
rect 1555 489 1579 506
rect 1555 472 1559 489
rect 1576 472 1579 489
rect 1555 455 1579 472
rect 1555 438 1559 455
rect 1576 438 1579 455
rect 1555 421 1579 438
rect 1555 404 1559 421
rect 1576 404 1579 421
rect 1555 387 1579 404
rect 1555 370 1559 387
rect 1576 370 1579 387
rect 1555 353 1579 370
rect 1555 336 1559 353
rect 1576 336 1579 353
rect 1555 319 1579 336
rect 1555 302 1559 319
rect 1576 302 1579 319
rect 1555 285 1579 302
rect 1555 268 1559 285
rect 1576 268 1579 285
rect 1555 251 1579 268
rect 1555 234 1559 251
rect 1576 234 1579 251
rect 1555 217 1579 234
rect 1555 200 1559 217
rect 1576 200 1579 217
rect 1555 183 1579 200
rect 1555 166 1559 183
rect 1576 166 1579 183
rect 1555 158 1579 166
rect 1600 1135 1624 1143
rect 1600 1118 1603 1135
rect 1620 1118 1624 1135
rect 1600 1101 1624 1118
rect 1600 1084 1603 1101
rect 1620 1084 1624 1101
rect 1600 1067 1624 1084
rect 1600 1050 1603 1067
rect 1620 1050 1624 1067
rect 1600 1033 1624 1050
rect 1600 1016 1603 1033
rect 1620 1016 1624 1033
rect 1600 999 1624 1016
rect 1600 982 1604 999
rect 1621 982 1624 999
rect 1600 965 1624 982
rect 1600 948 1604 965
rect 1621 948 1624 965
rect 1600 931 1624 948
rect 1600 914 1604 931
rect 1621 914 1624 931
rect 1600 897 1624 914
rect 1600 880 1604 897
rect 1621 880 1624 897
rect 1600 863 1624 880
rect 1600 846 1604 863
rect 1621 846 1624 863
rect 1600 829 1624 846
rect 1600 812 1604 829
rect 1621 812 1624 829
rect 1600 795 1624 812
rect 1600 778 1604 795
rect 1621 778 1624 795
rect 1600 761 1624 778
rect 1600 744 1604 761
rect 1621 744 1624 761
rect 1600 727 1624 744
rect 1600 710 1604 727
rect 1621 710 1624 727
rect 1600 693 1624 710
rect 1600 676 1604 693
rect 1621 676 1624 693
rect 1600 659 1624 676
rect 1600 642 1604 659
rect 1621 642 1624 659
rect 1600 625 1624 642
rect 1600 608 1604 625
rect 1621 608 1624 625
rect 1600 591 1624 608
rect 1600 574 1604 591
rect 1621 574 1624 591
rect 1600 557 1624 574
rect 1600 540 1604 557
rect 1621 540 1624 557
rect 1600 523 1624 540
rect 1600 506 1604 523
rect 1621 506 1624 523
rect 1600 489 1624 506
rect 1600 472 1604 489
rect 1621 472 1624 489
rect 1600 455 1624 472
rect 1600 438 1604 455
rect 1621 438 1624 455
rect 1600 421 1624 438
rect 1600 404 1604 421
rect 1621 404 1624 421
rect 1600 387 1624 404
rect 1600 370 1604 387
rect 1621 370 1624 387
rect 1600 353 1624 370
rect 1600 336 1604 353
rect 1621 336 1624 353
rect 1600 319 1624 336
rect 1600 302 1604 319
rect 1621 302 1624 319
rect 1600 285 1624 302
rect 1600 268 1604 285
rect 1621 268 1624 285
rect 1600 251 1624 268
rect 1600 234 1604 251
rect 1621 234 1624 251
rect 1600 217 1624 234
rect 1600 200 1604 217
rect 1621 200 1624 217
rect 1600 183 1624 200
rect 1600 166 1604 183
rect 1621 166 1624 183
rect 1600 115 1624 166
rect 1645 1135 1669 1184
rect 1645 1118 1648 1135
rect 1665 1118 1669 1135
rect 1645 1101 1669 1118
rect 1645 1084 1648 1101
rect 1665 1084 1669 1101
rect 1645 1067 1669 1084
rect 1645 1050 1648 1067
rect 1665 1050 1669 1067
rect 1645 1033 1669 1050
rect 1645 1016 1648 1033
rect 1665 1016 1669 1033
rect 1645 999 1669 1016
rect 1645 982 1649 999
rect 1666 982 1669 999
rect 1645 965 1669 982
rect 1645 948 1649 965
rect 1666 948 1669 965
rect 1645 931 1669 948
rect 1645 914 1649 931
rect 1666 914 1669 931
rect 1645 897 1669 914
rect 1645 880 1649 897
rect 1666 880 1669 897
rect 1645 863 1669 880
rect 1645 846 1649 863
rect 1666 846 1669 863
rect 1645 829 1669 846
rect 1645 812 1649 829
rect 1666 812 1669 829
rect 1645 795 1669 812
rect 1645 778 1649 795
rect 1666 778 1669 795
rect 1645 761 1669 778
rect 1645 744 1649 761
rect 1666 744 1669 761
rect 1645 727 1669 744
rect 1645 710 1649 727
rect 1666 710 1669 727
rect 1645 693 1669 710
rect 1645 676 1649 693
rect 1666 676 1669 693
rect 1645 659 1669 676
rect 1645 642 1649 659
rect 1666 642 1669 659
rect 1645 625 1669 642
rect 1645 608 1649 625
rect 1666 608 1669 625
rect 1645 591 1669 608
rect 1645 574 1649 591
rect 1666 574 1669 591
rect 1645 557 1669 574
rect 1645 540 1649 557
rect 1666 540 1669 557
rect 1645 523 1669 540
rect 1645 506 1649 523
rect 1666 506 1669 523
rect 1645 489 1669 506
rect 1645 472 1649 489
rect 1666 472 1669 489
rect 1645 455 1669 472
rect 1645 438 1649 455
rect 1666 438 1669 455
rect 1645 421 1669 438
rect 1645 404 1649 421
rect 1666 404 1669 421
rect 1645 387 1669 404
rect 1645 370 1649 387
rect 1666 370 1669 387
rect 1645 353 1669 370
rect 1645 336 1649 353
rect 1666 336 1669 353
rect 1645 319 1669 336
rect 1645 302 1649 319
rect 1666 302 1669 319
rect 1645 285 1669 302
rect 1645 268 1649 285
rect 1666 268 1669 285
rect 1645 251 1669 268
rect 1645 234 1649 251
rect 1666 234 1669 251
rect 1645 217 1669 234
rect 1645 200 1649 217
rect 1666 200 1669 217
rect 1645 183 1669 200
rect 1645 166 1649 183
rect 1666 166 1669 183
rect 1645 158 1669 166
rect 1690 1135 1714 1143
rect 1690 1118 1693 1135
rect 1710 1118 1714 1135
rect 1690 1101 1714 1118
rect 1690 1084 1693 1101
rect 1710 1084 1714 1101
rect 1690 1067 1714 1084
rect 1690 1050 1693 1067
rect 1710 1050 1714 1067
rect 1690 1033 1714 1050
rect 1690 1016 1693 1033
rect 1710 1016 1714 1033
rect 1690 999 1714 1016
rect 1690 982 1694 999
rect 1711 982 1714 999
rect 1690 965 1714 982
rect 1690 948 1694 965
rect 1711 948 1714 965
rect 1690 931 1714 948
rect 1690 914 1694 931
rect 1711 914 1714 931
rect 1690 897 1714 914
rect 1690 880 1694 897
rect 1711 880 1714 897
rect 1690 863 1714 880
rect 1690 846 1694 863
rect 1711 846 1714 863
rect 1690 829 1714 846
rect 1690 812 1694 829
rect 1711 812 1714 829
rect 1690 795 1714 812
rect 1690 778 1694 795
rect 1711 778 1714 795
rect 1690 761 1714 778
rect 1690 744 1694 761
rect 1711 744 1714 761
rect 1690 727 1714 744
rect 1690 710 1694 727
rect 1711 710 1714 727
rect 1690 693 1714 710
rect 1690 676 1694 693
rect 1711 676 1714 693
rect 1690 659 1714 676
rect 1690 642 1694 659
rect 1711 642 1714 659
rect 1690 625 1714 642
rect 1690 608 1694 625
rect 1711 608 1714 625
rect 1690 591 1714 608
rect 1690 574 1694 591
rect 1711 574 1714 591
rect 1690 557 1714 574
rect 1690 540 1694 557
rect 1711 540 1714 557
rect 1690 523 1714 540
rect 1690 506 1694 523
rect 1711 506 1714 523
rect 1690 489 1714 506
rect 1690 472 1694 489
rect 1711 472 1714 489
rect 1690 455 1714 472
rect 1690 438 1694 455
rect 1711 438 1714 455
rect 1690 421 1714 438
rect 1690 404 1694 421
rect 1711 404 1714 421
rect 1690 387 1714 404
rect 1690 370 1694 387
rect 1711 370 1714 387
rect 1690 353 1714 370
rect 1690 336 1694 353
rect 1711 336 1714 353
rect 1690 319 1714 336
rect 1690 302 1694 319
rect 1711 302 1714 319
rect 1690 285 1714 302
rect 1690 268 1694 285
rect 1711 268 1714 285
rect 1690 251 1714 268
rect 1690 234 1694 251
rect 1711 234 1714 251
rect 1690 217 1714 234
rect 1690 200 1694 217
rect 1711 200 1714 217
rect 1690 183 1714 200
rect 1690 166 1694 183
rect 1711 166 1714 183
rect 1690 115 1714 166
rect 1736 1135 1760 1184
rect 1736 1118 1739 1135
rect 1756 1118 1760 1135
rect 1736 1101 1760 1118
rect 1736 1084 1739 1101
rect 1756 1084 1760 1101
rect 1736 1067 1760 1084
rect 1736 1050 1739 1067
rect 1756 1050 1760 1067
rect 1736 1033 1760 1050
rect 1736 1016 1739 1033
rect 1756 1016 1760 1033
rect 1736 999 1760 1016
rect 1736 982 1740 999
rect 1757 982 1760 999
rect 1736 965 1760 982
rect 1736 948 1740 965
rect 1757 948 1760 965
rect 1736 931 1760 948
rect 1736 914 1740 931
rect 1757 914 1760 931
rect 1736 897 1760 914
rect 1736 880 1740 897
rect 1757 880 1760 897
rect 1736 863 1760 880
rect 1736 846 1740 863
rect 1757 846 1760 863
rect 1736 829 1760 846
rect 1736 812 1740 829
rect 1757 812 1760 829
rect 1736 795 1760 812
rect 1736 778 1740 795
rect 1757 778 1760 795
rect 1736 761 1760 778
rect 1736 744 1740 761
rect 1757 744 1760 761
rect 1736 727 1760 744
rect 1736 710 1740 727
rect 1757 710 1760 727
rect 1736 693 1760 710
rect 1736 676 1740 693
rect 1757 676 1760 693
rect 1736 659 1760 676
rect 1736 642 1740 659
rect 1757 642 1760 659
rect 1736 625 1760 642
rect 1736 608 1740 625
rect 1757 608 1760 625
rect 1736 591 1760 608
rect 1736 574 1740 591
rect 1757 574 1760 591
rect 1736 557 1760 574
rect 1736 540 1740 557
rect 1757 540 1760 557
rect 1736 523 1760 540
rect 1736 506 1740 523
rect 1757 506 1760 523
rect 1736 489 1760 506
rect 1736 472 1740 489
rect 1757 472 1760 489
rect 1736 455 1760 472
rect 1736 438 1740 455
rect 1757 438 1760 455
rect 1736 421 1760 438
rect 1736 404 1740 421
rect 1757 404 1760 421
rect 1736 387 1760 404
rect 1736 370 1740 387
rect 1757 370 1760 387
rect 1736 353 1760 370
rect 1736 336 1740 353
rect 1757 336 1760 353
rect 1736 319 1760 336
rect 1736 302 1740 319
rect 1757 302 1760 319
rect 1736 285 1760 302
rect 1736 268 1740 285
rect 1757 268 1760 285
rect 1736 251 1760 268
rect 1736 234 1740 251
rect 1757 234 1760 251
rect 1736 217 1760 234
rect 1736 200 1740 217
rect 1757 200 1760 217
rect 1736 183 1760 200
rect 1736 166 1740 183
rect 1757 166 1760 183
rect 1736 158 1760 166
rect 1781 1137 1804 1145
rect 1781 1120 1784 1137
rect 1801 1120 1804 1137
rect 1781 1103 1804 1120
rect 1781 1086 1784 1103
rect 1801 1086 1804 1103
rect 1781 1069 1804 1086
rect 1781 1052 1784 1069
rect 1801 1052 1804 1069
rect 1781 1035 1804 1052
rect 1781 1018 1784 1035
rect 1801 1018 1804 1035
rect 1781 1001 1804 1018
rect 1781 984 1784 1001
rect 1801 984 1804 1001
rect 1781 967 1804 984
rect 1781 950 1784 967
rect 1801 950 1804 967
rect 1781 933 1804 950
rect 1781 916 1784 933
rect 1801 916 1804 933
rect 1781 899 1804 916
rect 1781 882 1784 899
rect 1801 882 1804 899
rect 1781 865 1804 882
rect 1781 848 1784 865
rect 1801 848 1804 865
rect 1781 831 1804 848
rect 1781 814 1784 831
rect 1801 814 1804 831
rect 1781 797 1804 814
rect 1781 780 1784 797
rect 1801 780 1804 797
rect 1781 763 1804 780
rect 1781 746 1784 763
rect 1801 746 1804 763
rect 1781 729 1804 746
rect 1781 712 1784 729
rect 1801 712 1804 729
rect 1781 695 1804 712
rect 1781 678 1784 695
rect 1801 678 1804 695
rect 1781 661 1804 678
rect 1781 644 1784 661
rect 1801 644 1804 661
rect 1781 627 1804 644
rect 1781 610 1784 627
rect 1801 610 1804 627
rect 1781 593 1804 610
rect 1781 576 1784 593
rect 1801 576 1804 593
rect 1781 559 1804 576
rect 1781 542 1784 559
rect 1801 542 1804 559
rect 1781 525 1804 542
rect 1781 508 1784 525
rect 1801 508 1804 525
rect 1781 491 1804 508
rect 1781 474 1784 491
rect 1801 474 1804 491
rect 1781 457 1804 474
rect 1781 440 1784 457
rect 1801 440 1804 457
rect 1781 423 1804 440
rect 1781 406 1784 423
rect 1801 406 1804 423
rect 1781 389 1804 406
rect 1781 372 1784 389
rect 1801 372 1804 389
rect 1781 355 1804 372
rect 1781 338 1784 355
rect 1801 338 1804 355
rect 1781 321 1804 338
rect 1781 304 1784 321
rect 1801 304 1804 321
rect 1781 287 1804 304
rect 1781 270 1784 287
rect 1801 270 1804 287
rect 1781 253 1804 270
rect 1781 236 1784 253
rect 1801 236 1804 253
rect 1781 219 1804 236
rect 1781 202 1784 219
rect 1801 202 1804 219
rect 1781 185 1804 202
rect 1781 168 1784 185
rect 1801 168 1804 185
rect 1781 115 1804 168
rect 1825 1135 1849 1184
rect 1825 1118 1828 1135
rect 1845 1118 1849 1135
rect 1825 1101 1849 1118
rect 1825 1084 1828 1101
rect 1845 1084 1849 1101
rect 1825 1067 1849 1084
rect 1825 1050 1828 1067
rect 1845 1050 1849 1067
rect 1825 1033 1849 1050
rect 1825 1016 1828 1033
rect 1845 1016 1849 1033
rect 1825 999 1849 1016
rect 1825 982 1829 999
rect 1846 982 1849 999
rect 1825 965 1849 982
rect 1825 948 1829 965
rect 1846 948 1849 965
rect 1825 931 1849 948
rect 1825 914 1829 931
rect 1846 914 1849 931
rect 1825 897 1849 914
rect 1825 880 1829 897
rect 1846 880 1849 897
rect 1825 863 1849 880
rect 1825 846 1829 863
rect 1846 846 1849 863
rect 1825 829 1849 846
rect 1825 812 1829 829
rect 1846 812 1849 829
rect 1825 795 1849 812
rect 1825 778 1829 795
rect 1846 778 1849 795
rect 1825 761 1849 778
rect 1825 744 1829 761
rect 1846 744 1849 761
rect 1825 727 1849 744
rect 1825 710 1829 727
rect 1846 710 1849 727
rect 1825 693 1849 710
rect 1825 676 1829 693
rect 1846 676 1849 693
rect 1825 659 1849 676
rect 1825 642 1829 659
rect 1846 642 1849 659
rect 1825 625 1849 642
rect 1825 608 1829 625
rect 1846 608 1849 625
rect 1825 591 1849 608
rect 1825 574 1829 591
rect 1846 574 1849 591
rect 1825 557 1849 574
rect 1825 540 1829 557
rect 1846 540 1849 557
rect 1825 523 1849 540
rect 1825 506 1829 523
rect 1846 506 1849 523
rect 1825 489 1849 506
rect 1825 472 1829 489
rect 1846 472 1849 489
rect 1825 455 1849 472
rect 1825 438 1829 455
rect 1846 438 1849 455
rect 1825 421 1849 438
rect 1825 404 1829 421
rect 1846 404 1849 421
rect 1825 387 1849 404
rect 1825 370 1829 387
rect 1846 370 1849 387
rect 1825 353 1849 370
rect 1825 336 1829 353
rect 1846 336 1849 353
rect 1825 319 1849 336
rect 1825 302 1829 319
rect 1846 302 1849 319
rect 1825 285 1849 302
rect 1825 268 1829 285
rect 1846 268 1849 285
rect 1825 251 1849 268
rect 1825 234 1829 251
rect 1846 234 1849 251
rect 1825 217 1849 234
rect 1825 200 1829 217
rect 1846 200 1849 217
rect 1825 183 1849 200
rect 1825 166 1829 183
rect 1846 166 1849 183
rect 1825 158 1849 166
rect 1870 1135 1894 1143
rect 1870 1118 1873 1135
rect 1890 1118 1894 1135
rect 1870 1101 1894 1118
rect 1870 1084 1873 1101
rect 1890 1084 1894 1101
rect 1870 1067 1894 1084
rect 1870 1050 1873 1067
rect 1890 1050 1894 1067
rect 1870 1033 1894 1050
rect 1870 1016 1873 1033
rect 1890 1016 1894 1033
rect 1870 999 1894 1016
rect 1870 982 1874 999
rect 1891 982 1894 999
rect 1870 965 1894 982
rect 1870 948 1874 965
rect 1891 948 1894 965
rect 1870 931 1894 948
rect 1870 914 1874 931
rect 1891 914 1894 931
rect 1870 897 1894 914
rect 1870 880 1874 897
rect 1891 880 1894 897
rect 1870 863 1894 880
rect 1870 846 1874 863
rect 1891 846 1894 863
rect 1870 829 1894 846
rect 1870 812 1874 829
rect 1891 812 1894 829
rect 1870 795 1894 812
rect 1870 778 1874 795
rect 1891 778 1894 795
rect 1870 761 1894 778
rect 1870 744 1874 761
rect 1891 744 1894 761
rect 1870 727 1894 744
rect 1870 710 1874 727
rect 1891 710 1894 727
rect 1870 693 1894 710
rect 1870 676 1874 693
rect 1891 676 1894 693
rect 1870 659 1894 676
rect 1870 642 1874 659
rect 1891 642 1894 659
rect 1870 625 1894 642
rect 1870 608 1874 625
rect 1891 608 1894 625
rect 1870 591 1894 608
rect 1870 574 1874 591
rect 1891 574 1894 591
rect 1870 557 1894 574
rect 1870 540 1874 557
rect 1891 540 1894 557
rect 1870 523 1894 540
rect 1870 506 1874 523
rect 1891 506 1894 523
rect 1870 489 1894 506
rect 1870 472 1874 489
rect 1891 472 1894 489
rect 1870 455 1894 472
rect 1870 438 1874 455
rect 1891 438 1894 455
rect 1870 421 1894 438
rect 1870 404 1874 421
rect 1891 404 1894 421
rect 1870 387 1894 404
rect 1870 370 1874 387
rect 1891 370 1894 387
rect 1870 353 1894 370
rect 1870 336 1874 353
rect 1891 336 1894 353
rect 1870 319 1894 336
rect 1870 302 1874 319
rect 1891 302 1894 319
rect 1870 285 1894 302
rect 1870 268 1874 285
rect 1891 268 1894 285
rect 1870 251 1894 268
rect 1870 234 1874 251
rect 1891 234 1894 251
rect 1870 217 1894 234
rect 1870 200 1874 217
rect 1891 200 1894 217
rect 1870 183 1894 200
rect 1870 166 1874 183
rect 1891 166 1894 183
rect 1870 115 1894 166
rect 1915 1135 1939 1184
rect 1915 1118 1918 1135
rect 1935 1118 1939 1135
rect 1915 1101 1939 1118
rect 1915 1084 1918 1101
rect 1935 1084 1939 1101
rect 1915 1067 1939 1084
rect 1915 1050 1918 1067
rect 1935 1050 1939 1067
rect 1915 1033 1939 1050
rect 1915 1016 1918 1033
rect 1935 1016 1939 1033
rect 1915 999 1939 1016
rect 1915 982 1919 999
rect 1936 982 1939 999
rect 1915 965 1939 982
rect 1915 948 1919 965
rect 1936 948 1939 965
rect 1915 931 1939 948
rect 1915 914 1919 931
rect 1936 914 1939 931
rect 1915 897 1939 914
rect 1915 880 1919 897
rect 1936 880 1939 897
rect 1915 863 1939 880
rect 1915 846 1919 863
rect 1936 846 1939 863
rect 1915 829 1939 846
rect 1915 812 1919 829
rect 1936 812 1939 829
rect 1915 795 1939 812
rect 1915 778 1919 795
rect 1936 778 1939 795
rect 1915 761 1939 778
rect 1915 744 1919 761
rect 1936 744 1939 761
rect 1915 727 1939 744
rect 1915 710 1919 727
rect 1936 710 1939 727
rect 1915 693 1939 710
rect 1915 676 1919 693
rect 1936 676 1939 693
rect 1915 659 1939 676
rect 1915 642 1919 659
rect 1936 642 1939 659
rect 1915 625 1939 642
rect 1915 608 1919 625
rect 1936 608 1939 625
rect 1915 591 1939 608
rect 1915 574 1919 591
rect 1936 574 1939 591
rect 1915 557 1939 574
rect 1915 540 1919 557
rect 1936 540 1939 557
rect 1915 523 1939 540
rect 1915 506 1919 523
rect 1936 506 1939 523
rect 1915 489 1939 506
rect 1915 472 1919 489
rect 1936 472 1939 489
rect 1915 455 1939 472
rect 1915 438 1919 455
rect 1936 438 1939 455
rect 1915 421 1939 438
rect 1915 404 1919 421
rect 1936 404 1939 421
rect 1915 387 1939 404
rect 1915 370 1919 387
rect 1936 370 1939 387
rect 1915 353 1939 370
rect 1915 336 1919 353
rect 1936 336 1939 353
rect 1915 319 1939 336
rect 1915 302 1919 319
rect 1936 302 1939 319
rect 1915 285 1939 302
rect 1915 268 1919 285
rect 1936 268 1939 285
rect 1915 251 1939 268
rect 1915 234 1919 251
rect 1936 234 1939 251
rect 1915 217 1939 234
rect 1915 200 1919 217
rect 1936 200 1939 217
rect 1915 183 1939 200
rect 1915 166 1919 183
rect 1936 166 1939 183
rect 1915 158 1939 166
rect 1960 1135 1984 1143
rect 1960 1118 1963 1135
rect 1980 1118 1984 1135
rect 1960 1101 1984 1118
rect 1960 1084 1963 1101
rect 1980 1084 1984 1101
rect 1960 1067 1984 1084
rect 1960 1050 1963 1067
rect 1980 1050 1984 1067
rect 1960 1033 1984 1050
rect 1960 1016 1963 1033
rect 1980 1016 1984 1033
rect 1960 999 1984 1016
rect 1960 982 1964 999
rect 1981 982 1984 999
rect 1960 965 1984 982
rect 1960 948 1964 965
rect 1981 948 1984 965
rect 1960 931 1984 948
rect 1960 914 1964 931
rect 1981 914 1984 931
rect 1960 897 1984 914
rect 1960 880 1964 897
rect 1981 880 1984 897
rect 1960 863 1984 880
rect 1960 846 1964 863
rect 1981 846 1984 863
rect 1960 829 1984 846
rect 1960 812 1964 829
rect 1981 812 1984 829
rect 1960 795 1984 812
rect 1960 778 1964 795
rect 1981 778 1984 795
rect 1960 761 1984 778
rect 1960 744 1964 761
rect 1981 744 1984 761
rect 1960 727 1984 744
rect 1960 710 1964 727
rect 1981 710 1984 727
rect 1960 693 1984 710
rect 1960 676 1964 693
rect 1981 676 1984 693
rect 1960 659 1984 676
rect 1960 642 1964 659
rect 1981 642 1984 659
rect 1960 625 1984 642
rect 1960 608 1964 625
rect 1981 608 1984 625
rect 1960 591 1984 608
rect 1960 574 1964 591
rect 1981 574 1984 591
rect 1960 557 1984 574
rect 1960 540 1964 557
rect 1981 540 1984 557
rect 1960 523 1984 540
rect 1960 506 1964 523
rect 1981 506 1984 523
rect 1960 489 1984 506
rect 1960 472 1964 489
rect 1981 472 1984 489
rect 1960 455 1984 472
rect 1960 438 1964 455
rect 1981 438 1984 455
rect 1960 421 1984 438
rect 1960 404 1964 421
rect 1981 404 1984 421
rect 1960 387 1984 404
rect 1960 370 1964 387
rect 1981 370 1984 387
rect 1960 353 1984 370
rect 1960 336 1964 353
rect 1981 336 1984 353
rect 1960 319 1984 336
rect 1960 302 1964 319
rect 1981 302 1984 319
rect 1960 285 1984 302
rect 1960 268 1964 285
rect 1981 268 1984 285
rect 1960 251 1984 268
rect 1960 234 1964 251
rect 1981 234 1984 251
rect 1960 217 1984 234
rect 1960 200 1964 217
rect 1981 200 1984 217
rect 1960 183 1984 200
rect 1960 166 1964 183
rect 1981 166 1984 183
rect 1960 115 1984 166
rect 2005 1135 2029 1184
rect 2005 1118 2008 1135
rect 2025 1118 2029 1135
rect 2005 1101 2029 1118
rect 2005 1084 2008 1101
rect 2025 1084 2029 1101
rect 2005 1067 2029 1084
rect 2005 1050 2008 1067
rect 2025 1050 2029 1067
rect 2005 1033 2029 1050
rect 2005 1016 2008 1033
rect 2025 1016 2029 1033
rect 2005 999 2029 1016
rect 2005 982 2009 999
rect 2026 982 2029 999
rect 2005 965 2029 982
rect 2005 948 2009 965
rect 2026 948 2029 965
rect 2005 931 2029 948
rect 2005 914 2009 931
rect 2026 914 2029 931
rect 2005 897 2029 914
rect 2005 880 2009 897
rect 2026 880 2029 897
rect 2005 863 2029 880
rect 2005 846 2009 863
rect 2026 846 2029 863
rect 2005 829 2029 846
rect 2005 812 2009 829
rect 2026 812 2029 829
rect 2005 795 2029 812
rect 2005 778 2009 795
rect 2026 778 2029 795
rect 2005 761 2029 778
rect 2005 744 2009 761
rect 2026 744 2029 761
rect 2005 727 2029 744
rect 2005 710 2009 727
rect 2026 710 2029 727
rect 2005 693 2029 710
rect 2005 676 2009 693
rect 2026 676 2029 693
rect 2005 659 2029 676
rect 2005 642 2009 659
rect 2026 642 2029 659
rect 2005 625 2029 642
rect 2005 608 2009 625
rect 2026 608 2029 625
rect 2005 591 2029 608
rect 2005 574 2009 591
rect 2026 574 2029 591
rect 2005 557 2029 574
rect 2005 540 2009 557
rect 2026 540 2029 557
rect 2005 523 2029 540
rect 2005 506 2009 523
rect 2026 506 2029 523
rect 2005 489 2029 506
rect 2005 472 2009 489
rect 2026 472 2029 489
rect 2005 455 2029 472
rect 2005 438 2009 455
rect 2026 438 2029 455
rect 2005 421 2029 438
rect 2005 404 2009 421
rect 2026 404 2029 421
rect 2005 387 2029 404
rect 2005 370 2009 387
rect 2026 370 2029 387
rect 2005 353 2029 370
rect 2005 336 2009 353
rect 2026 336 2029 353
rect 2005 319 2029 336
rect 2005 302 2009 319
rect 2026 302 2029 319
rect 2005 285 2029 302
rect 2005 268 2009 285
rect 2026 268 2029 285
rect 2005 251 2029 268
rect 2005 234 2009 251
rect 2026 234 2029 251
rect 2005 217 2029 234
rect 2005 200 2009 217
rect 2026 200 2029 217
rect 2005 183 2029 200
rect 2005 166 2009 183
rect 2026 166 2029 183
rect 2005 158 2029 166
rect 2050 1135 2074 1143
rect 2050 1118 2053 1135
rect 2070 1118 2074 1135
rect 2050 1101 2074 1118
rect 2050 1084 2053 1101
rect 2070 1084 2074 1101
rect 2050 1067 2074 1084
rect 2050 1050 2053 1067
rect 2070 1050 2074 1067
rect 2050 1033 2074 1050
rect 2050 1016 2053 1033
rect 2070 1016 2074 1033
rect 2050 999 2074 1016
rect 2050 982 2054 999
rect 2071 982 2074 999
rect 2050 965 2074 982
rect 2050 948 2054 965
rect 2071 948 2074 965
rect 2050 931 2074 948
rect 2050 914 2054 931
rect 2071 914 2074 931
rect 2050 897 2074 914
rect 2050 880 2054 897
rect 2071 880 2074 897
rect 2050 863 2074 880
rect 2050 846 2054 863
rect 2071 846 2074 863
rect 2050 829 2074 846
rect 2050 812 2054 829
rect 2071 812 2074 829
rect 2050 795 2074 812
rect 2050 778 2054 795
rect 2071 778 2074 795
rect 2050 761 2074 778
rect 2050 744 2054 761
rect 2071 744 2074 761
rect 2050 727 2074 744
rect 2050 710 2054 727
rect 2071 710 2074 727
rect 2050 693 2074 710
rect 2050 676 2054 693
rect 2071 676 2074 693
rect 2050 659 2074 676
rect 2050 642 2054 659
rect 2071 642 2074 659
rect 2050 625 2074 642
rect 2050 608 2054 625
rect 2071 608 2074 625
rect 2050 591 2074 608
rect 2050 574 2054 591
rect 2071 574 2074 591
rect 2050 557 2074 574
rect 2050 540 2054 557
rect 2071 540 2074 557
rect 2050 523 2074 540
rect 2050 506 2054 523
rect 2071 506 2074 523
rect 2050 489 2074 506
rect 2050 472 2054 489
rect 2071 472 2074 489
rect 2050 455 2074 472
rect 2050 438 2054 455
rect 2071 438 2074 455
rect 2050 421 2074 438
rect 2050 404 2054 421
rect 2071 404 2074 421
rect 2050 387 2074 404
rect 2050 370 2054 387
rect 2071 370 2074 387
rect 2050 353 2074 370
rect 2050 336 2054 353
rect 2071 336 2074 353
rect 2050 319 2074 336
rect 2050 302 2054 319
rect 2071 302 2074 319
rect 2050 285 2074 302
rect 2050 268 2054 285
rect 2071 268 2074 285
rect 2050 251 2074 268
rect 2050 234 2054 251
rect 2071 234 2074 251
rect 2050 217 2074 234
rect 2050 200 2054 217
rect 2071 200 2074 217
rect 2050 183 2074 200
rect 2050 166 2054 183
rect 2071 166 2074 183
rect 2050 115 2074 166
rect 2095 1135 2119 1184
rect 2095 1118 2098 1135
rect 2115 1118 2119 1135
rect 2095 1101 2119 1118
rect 2095 1084 2098 1101
rect 2115 1084 2119 1101
rect 2095 1067 2119 1084
rect 2095 1050 2098 1067
rect 2115 1050 2119 1067
rect 2095 1033 2119 1050
rect 2095 1016 2098 1033
rect 2115 1016 2119 1033
rect 2095 999 2119 1016
rect 2095 982 2099 999
rect 2116 982 2119 999
rect 2095 965 2119 982
rect 2095 948 2099 965
rect 2116 948 2119 965
rect 2095 931 2119 948
rect 2095 914 2099 931
rect 2116 914 2119 931
rect 2095 897 2119 914
rect 2095 880 2099 897
rect 2116 880 2119 897
rect 2095 863 2119 880
rect 2095 846 2099 863
rect 2116 846 2119 863
rect 2095 829 2119 846
rect 2095 812 2099 829
rect 2116 812 2119 829
rect 2095 795 2119 812
rect 2095 778 2099 795
rect 2116 778 2119 795
rect 2095 761 2119 778
rect 2095 744 2099 761
rect 2116 744 2119 761
rect 2095 727 2119 744
rect 2095 710 2099 727
rect 2116 710 2119 727
rect 2095 693 2119 710
rect 2095 676 2099 693
rect 2116 676 2119 693
rect 2095 659 2119 676
rect 2095 642 2099 659
rect 2116 642 2119 659
rect 2095 625 2119 642
rect 2095 608 2099 625
rect 2116 608 2119 625
rect 2095 591 2119 608
rect 2095 574 2099 591
rect 2116 574 2119 591
rect 2095 557 2119 574
rect 2095 540 2099 557
rect 2116 540 2119 557
rect 2095 523 2119 540
rect 2095 506 2099 523
rect 2116 506 2119 523
rect 2095 489 2119 506
rect 2095 472 2099 489
rect 2116 472 2119 489
rect 2095 455 2119 472
rect 2095 438 2099 455
rect 2116 438 2119 455
rect 2095 421 2119 438
rect 2095 404 2099 421
rect 2116 404 2119 421
rect 2095 387 2119 404
rect 2095 370 2099 387
rect 2116 370 2119 387
rect 2095 353 2119 370
rect 2095 336 2099 353
rect 2116 336 2119 353
rect 2095 319 2119 336
rect 2095 302 2099 319
rect 2116 302 2119 319
rect 2095 285 2119 302
rect 2095 268 2099 285
rect 2116 268 2119 285
rect 2095 251 2119 268
rect 2095 234 2099 251
rect 2116 234 2119 251
rect 2095 217 2119 234
rect 2095 200 2099 217
rect 2116 200 2119 217
rect 2095 183 2119 200
rect 2095 166 2099 183
rect 2116 166 2119 183
rect 2095 158 2119 166
rect 2140 1137 2163 1145
rect 2140 1120 2143 1137
rect 2160 1120 2163 1137
rect 2140 1103 2163 1120
rect 2140 1086 2143 1103
rect 2160 1086 2163 1103
rect 2140 1069 2163 1086
rect 2140 1052 2143 1069
rect 2160 1052 2163 1069
rect 2140 1035 2163 1052
rect 2140 1018 2143 1035
rect 2160 1018 2163 1035
rect 2140 1001 2163 1018
rect 2140 984 2143 1001
rect 2160 984 2163 1001
rect 2140 967 2163 984
rect 2140 950 2143 967
rect 2160 950 2163 967
rect 2140 933 2163 950
rect 2140 916 2143 933
rect 2160 916 2163 933
rect 2140 899 2163 916
rect 2140 882 2143 899
rect 2160 882 2163 899
rect 2140 865 2163 882
rect 2140 848 2143 865
rect 2160 848 2163 865
rect 2140 831 2163 848
rect 2140 814 2143 831
rect 2160 814 2163 831
rect 2140 797 2163 814
rect 2140 780 2143 797
rect 2160 780 2163 797
rect 2140 763 2163 780
rect 2140 746 2143 763
rect 2160 746 2163 763
rect 2140 729 2163 746
rect 2140 712 2143 729
rect 2160 712 2163 729
rect 2140 695 2163 712
rect 2140 678 2143 695
rect 2160 678 2163 695
rect 2140 661 2163 678
rect 2140 644 2143 661
rect 2160 644 2163 661
rect 2140 627 2163 644
rect 2140 610 2143 627
rect 2160 610 2163 627
rect 2140 593 2163 610
rect 2140 576 2143 593
rect 2160 576 2163 593
rect 2140 559 2163 576
rect 2140 542 2143 559
rect 2160 542 2163 559
rect 2140 525 2163 542
rect 2140 508 2143 525
rect 2160 508 2163 525
rect 2140 491 2163 508
rect 2140 474 2143 491
rect 2160 474 2163 491
rect 2140 457 2163 474
rect 2140 440 2143 457
rect 2160 440 2163 457
rect 2140 423 2163 440
rect 2140 406 2143 423
rect 2160 406 2163 423
rect 2140 389 2163 406
rect 2140 372 2143 389
rect 2160 372 2163 389
rect 2140 355 2163 372
rect 2140 338 2143 355
rect 2160 338 2163 355
rect 2140 321 2163 338
rect 2140 304 2143 321
rect 2160 304 2163 321
rect 2140 287 2163 304
rect 2140 270 2143 287
rect 2160 270 2163 287
rect 2140 253 2163 270
rect 2140 236 2143 253
rect 2160 236 2163 253
rect 2140 219 2163 236
rect 2140 202 2143 219
rect 2160 202 2163 219
rect 2140 185 2163 202
rect 2140 168 2143 185
rect 2160 168 2163 185
rect 2140 115 2163 168
rect 2184 1135 2208 1184
rect 2184 1118 2187 1135
rect 2204 1118 2208 1135
rect 2184 1101 2208 1118
rect 2184 1084 2187 1101
rect 2204 1084 2208 1101
rect 2184 1067 2208 1084
rect 2184 1050 2187 1067
rect 2204 1050 2208 1067
rect 2184 1033 2208 1050
rect 2184 1016 2187 1033
rect 2204 1016 2208 1033
rect 2184 999 2208 1016
rect 2184 982 2188 999
rect 2205 982 2208 999
rect 2184 965 2208 982
rect 2184 948 2188 965
rect 2205 948 2208 965
rect 2184 931 2208 948
rect 2184 914 2188 931
rect 2205 914 2208 931
rect 2184 897 2208 914
rect 2184 880 2188 897
rect 2205 880 2208 897
rect 2184 863 2208 880
rect 2184 846 2188 863
rect 2205 846 2208 863
rect 2184 829 2208 846
rect 2184 812 2188 829
rect 2205 812 2208 829
rect 2184 795 2208 812
rect 2184 778 2188 795
rect 2205 778 2208 795
rect 2184 761 2208 778
rect 2184 744 2188 761
rect 2205 744 2208 761
rect 2184 727 2208 744
rect 2184 710 2188 727
rect 2205 710 2208 727
rect 2184 693 2208 710
rect 2184 676 2188 693
rect 2205 676 2208 693
rect 2184 659 2208 676
rect 2184 642 2188 659
rect 2205 642 2208 659
rect 2184 625 2208 642
rect 2184 608 2188 625
rect 2205 608 2208 625
rect 2184 591 2208 608
rect 2184 574 2188 591
rect 2205 574 2208 591
rect 2184 557 2208 574
rect 2184 540 2188 557
rect 2205 540 2208 557
rect 2184 523 2208 540
rect 2184 506 2188 523
rect 2205 506 2208 523
rect 2184 489 2208 506
rect 2184 472 2188 489
rect 2205 472 2208 489
rect 2184 455 2208 472
rect 2184 438 2188 455
rect 2205 438 2208 455
rect 2184 421 2208 438
rect 2184 404 2188 421
rect 2205 404 2208 421
rect 2184 387 2208 404
rect 2184 370 2188 387
rect 2205 370 2208 387
rect 2184 353 2208 370
rect 2184 336 2188 353
rect 2205 336 2208 353
rect 2184 319 2208 336
rect 2184 302 2188 319
rect 2205 302 2208 319
rect 2184 285 2208 302
rect 2184 268 2188 285
rect 2205 268 2208 285
rect 2184 251 2208 268
rect 2184 234 2188 251
rect 2205 234 2208 251
rect 2184 217 2208 234
rect 2184 200 2188 217
rect 2205 200 2208 217
rect 2184 183 2208 200
rect 2184 166 2188 183
rect 2205 166 2208 183
rect 2184 158 2208 166
rect 2229 1135 2253 1143
rect 2229 1118 2232 1135
rect 2249 1118 2253 1135
rect 2229 1101 2253 1118
rect 2229 1084 2232 1101
rect 2249 1084 2253 1101
rect 2229 1067 2253 1084
rect 2229 1050 2232 1067
rect 2249 1050 2253 1067
rect 2229 1033 2253 1050
rect 2229 1016 2232 1033
rect 2249 1016 2253 1033
rect 2229 999 2253 1016
rect 2229 982 2233 999
rect 2250 982 2253 999
rect 2229 965 2253 982
rect 2229 948 2233 965
rect 2250 948 2253 965
rect 2229 931 2253 948
rect 2229 914 2233 931
rect 2250 914 2253 931
rect 2229 897 2253 914
rect 2229 880 2233 897
rect 2250 880 2253 897
rect 2229 863 2253 880
rect 2229 846 2233 863
rect 2250 846 2253 863
rect 2229 829 2253 846
rect 2229 812 2233 829
rect 2250 812 2253 829
rect 2229 795 2253 812
rect 2229 778 2233 795
rect 2250 778 2253 795
rect 2229 761 2253 778
rect 2229 744 2233 761
rect 2250 744 2253 761
rect 2229 727 2253 744
rect 2229 710 2233 727
rect 2250 710 2253 727
rect 2229 693 2253 710
rect 2229 676 2233 693
rect 2250 676 2253 693
rect 2229 659 2253 676
rect 2229 642 2233 659
rect 2250 642 2253 659
rect 2229 625 2253 642
rect 2229 608 2233 625
rect 2250 608 2253 625
rect 2229 591 2253 608
rect 2229 574 2233 591
rect 2250 574 2253 591
rect 2229 557 2253 574
rect 2229 540 2233 557
rect 2250 540 2253 557
rect 2229 523 2253 540
rect 2229 506 2233 523
rect 2250 506 2253 523
rect 2229 489 2253 506
rect 2229 472 2233 489
rect 2250 472 2253 489
rect 2229 455 2253 472
rect 2229 438 2233 455
rect 2250 438 2253 455
rect 2229 421 2253 438
rect 2229 404 2233 421
rect 2250 404 2253 421
rect 2229 387 2253 404
rect 2229 370 2233 387
rect 2250 370 2253 387
rect 2229 353 2253 370
rect 2229 336 2233 353
rect 2250 336 2253 353
rect 2229 319 2253 336
rect 2229 302 2233 319
rect 2250 302 2253 319
rect 2229 285 2253 302
rect 2229 268 2233 285
rect 2250 268 2253 285
rect 2229 251 2253 268
rect 2229 234 2233 251
rect 2250 234 2253 251
rect 2229 217 2253 234
rect 2229 200 2233 217
rect 2250 200 2253 217
rect 2229 183 2253 200
rect 2229 166 2233 183
rect 2250 166 2253 183
rect 2229 115 2253 166
rect 2274 1135 2298 1184
rect 2274 1118 2277 1135
rect 2294 1118 2298 1135
rect 2274 1101 2298 1118
rect 2274 1084 2277 1101
rect 2294 1084 2298 1101
rect 2274 1067 2298 1084
rect 2274 1050 2277 1067
rect 2294 1050 2298 1067
rect 2274 1033 2298 1050
rect 2274 1016 2277 1033
rect 2294 1016 2298 1033
rect 2274 999 2298 1016
rect 2274 982 2278 999
rect 2295 982 2298 999
rect 2274 965 2298 982
rect 2274 948 2278 965
rect 2295 948 2298 965
rect 2274 931 2298 948
rect 2274 914 2278 931
rect 2295 914 2298 931
rect 2274 897 2298 914
rect 2274 880 2278 897
rect 2295 880 2298 897
rect 2274 863 2298 880
rect 2274 846 2278 863
rect 2295 846 2298 863
rect 2274 829 2298 846
rect 2274 812 2278 829
rect 2295 812 2298 829
rect 2274 795 2298 812
rect 2274 778 2278 795
rect 2295 778 2298 795
rect 2274 761 2298 778
rect 2274 744 2278 761
rect 2295 744 2298 761
rect 2274 727 2298 744
rect 2274 710 2278 727
rect 2295 710 2298 727
rect 2274 693 2298 710
rect 2274 676 2278 693
rect 2295 676 2298 693
rect 2274 659 2298 676
rect 2274 642 2278 659
rect 2295 642 2298 659
rect 2274 625 2298 642
rect 2274 608 2278 625
rect 2295 608 2298 625
rect 2274 591 2298 608
rect 2274 574 2278 591
rect 2295 574 2298 591
rect 2274 557 2298 574
rect 2274 540 2278 557
rect 2295 540 2298 557
rect 2274 523 2298 540
rect 2274 506 2278 523
rect 2295 506 2298 523
rect 2274 489 2298 506
rect 2274 472 2278 489
rect 2295 472 2298 489
rect 2274 455 2298 472
rect 2274 438 2278 455
rect 2295 438 2298 455
rect 2274 421 2298 438
rect 2274 404 2278 421
rect 2295 404 2298 421
rect 2274 387 2298 404
rect 2274 370 2278 387
rect 2295 370 2298 387
rect 2274 353 2298 370
rect 2274 336 2278 353
rect 2295 336 2298 353
rect 2274 319 2298 336
rect 2274 302 2278 319
rect 2295 302 2298 319
rect 2274 285 2298 302
rect 2274 268 2278 285
rect 2295 268 2298 285
rect 2274 251 2298 268
rect 2274 234 2278 251
rect 2295 234 2298 251
rect 2274 217 2298 234
rect 2274 200 2278 217
rect 2295 200 2298 217
rect 2274 183 2298 200
rect 2274 166 2278 183
rect 2295 166 2298 183
rect 2274 158 2298 166
rect 2319 1135 2343 1143
rect 2319 1118 2322 1135
rect 2339 1118 2343 1135
rect 2319 1101 2343 1118
rect 2319 1084 2322 1101
rect 2339 1084 2343 1101
rect 2319 1067 2343 1084
rect 2319 1050 2322 1067
rect 2339 1050 2343 1067
rect 2319 1033 2343 1050
rect 2319 1016 2322 1033
rect 2339 1016 2343 1033
rect 2319 999 2343 1016
rect 2319 982 2323 999
rect 2340 982 2343 999
rect 2319 965 2343 982
rect 2319 948 2323 965
rect 2340 948 2343 965
rect 2319 931 2343 948
rect 2319 914 2323 931
rect 2340 914 2343 931
rect 2319 897 2343 914
rect 2319 880 2323 897
rect 2340 880 2343 897
rect 2319 863 2343 880
rect 2319 846 2323 863
rect 2340 846 2343 863
rect 2319 829 2343 846
rect 2319 812 2323 829
rect 2340 812 2343 829
rect 2319 795 2343 812
rect 2319 778 2323 795
rect 2340 778 2343 795
rect 2319 761 2343 778
rect 2319 744 2323 761
rect 2340 744 2343 761
rect 2319 727 2343 744
rect 2319 710 2323 727
rect 2340 710 2343 727
rect 2319 693 2343 710
rect 2319 676 2323 693
rect 2340 676 2343 693
rect 2319 659 2343 676
rect 2319 642 2323 659
rect 2340 642 2343 659
rect 2319 625 2343 642
rect 2319 608 2323 625
rect 2340 608 2343 625
rect 2319 591 2343 608
rect 2319 574 2323 591
rect 2340 574 2343 591
rect 2319 557 2343 574
rect 2319 540 2323 557
rect 2340 540 2343 557
rect 2319 523 2343 540
rect 2319 506 2323 523
rect 2340 506 2343 523
rect 2319 489 2343 506
rect 2319 472 2323 489
rect 2340 472 2343 489
rect 2319 455 2343 472
rect 2319 438 2323 455
rect 2340 438 2343 455
rect 2319 421 2343 438
rect 2319 404 2323 421
rect 2340 404 2343 421
rect 2319 387 2343 404
rect 2319 370 2323 387
rect 2340 370 2343 387
rect 2319 353 2343 370
rect 2319 336 2323 353
rect 2340 336 2343 353
rect 2319 319 2343 336
rect 2319 302 2323 319
rect 2340 302 2343 319
rect 2319 285 2343 302
rect 2319 268 2323 285
rect 2340 268 2343 285
rect 2319 251 2343 268
rect 2319 234 2323 251
rect 2340 234 2343 251
rect 2319 217 2343 234
rect 2319 200 2323 217
rect 2340 200 2343 217
rect 2319 183 2343 200
rect 2319 166 2323 183
rect 2340 166 2343 183
rect 2319 115 2343 166
rect 2364 1135 2388 1184
rect 2364 1118 2367 1135
rect 2384 1118 2388 1135
rect 2364 1101 2388 1118
rect 2364 1084 2367 1101
rect 2384 1084 2388 1101
rect 2364 1067 2388 1084
rect 2364 1050 2367 1067
rect 2384 1050 2388 1067
rect 2364 1033 2388 1050
rect 2364 1016 2367 1033
rect 2384 1016 2388 1033
rect 2364 999 2388 1016
rect 2364 982 2368 999
rect 2385 982 2388 999
rect 2364 965 2388 982
rect 2364 948 2368 965
rect 2385 948 2388 965
rect 2364 931 2388 948
rect 2364 914 2368 931
rect 2385 914 2388 931
rect 2364 897 2388 914
rect 2364 880 2368 897
rect 2385 880 2388 897
rect 2364 863 2388 880
rect 2364 846 2368 863
rect 2385 846 2388 863
rect 2364 829 2388 846
rect 2364 812 2368 829
rect 2385 812 2388 829
rect 2364 795 2388 812
rect 2364 778 2368 795
rect 2385 778 2388 795
rect 2364 761 2388 778
rect 2364 744 2368 761
rect 2385 744 2388 761
rect 2364 727 2388 744
rect 2364 710 2368 727
rect 2385 710 2388 727
rect 2364 693 2388 710
rect 2364 676 2368 693
rect 2385 676 2388 693
rect 2364 659 2388 676
rect 2364 642 2368 659
rect 2385 642 2388 659
rect 2364 625 2388 642
rect 2364 608 2368 625
rect 2385 608 2388 625
rect 2364 591 2388 608
rect 2364 574 2368 591
rect 2385 574 2388 591
rect 2364 557 2388 574
rect 2364 540 2368 557
rect 2385 540 2388 557
rect 2364 523 2388 540
rect 2364 506 2368 523
rect 2385 506 2388 523
rect 2364 489 2388 506
rect 2364 472 2368 489
rect 2385 472 2388 489
rect 2364 455 2388 472
rect 2364 438 2368 455
rect 2385 438 2388 455
rect 2364 421 2388 438
rect 2364 404 2368 421
rect 2385 404 2388 421
rect 2364 387 2388 404
rect 2364 370 2368 387
rect 2385 370 2388 387
rect 2364 353 2388 370
rect 2364 336 2368 353
rect 2385 336 2388 353
rect 2364 319 2388 336
rect 2364 302 2368 319
rect 2385 302 2388 319
rect 2364 285 2388 302
rect 2364 268 2368 285
rect 2385 268 2388 285
rect 2364 251 2388 268
rect 2364 234 2368 251
rect 2385 234 2388 251
rect 2364 217 2388 234
rect 2364 200 2368 217
rect 2385 200 2388 217
rect 2364 183 2388 200
rect 2364 166 2368 183
rect 2385 166 2388 183
rect 2364 158 2388 166
rect 2409 1135 2433 1143
rect 2409 1118 2412 1135
rect 2429 1118 2433 1135
rect 2409 1101 2433 1118
rect 2409 1084 2412 1101
rect 2429 1084 2433 1101
rect 2409 1067 2433 1084
rect 2409 1050 2412 1067
rect 2429 1050 2433 1067
rect 2409 1033 2433 1050
rect 2409 1016 2412 1033
rect 2429 1016 2433 1033
rect 2409 999 2433 1016
rect 2409 982 2413 999
rect 2430 982 2433 999
rect 2409 965 2433 982
rect 2409 948 2413 965
rect 2430 948 2433 965
rect 2409 931 2433 948
rect 2409 914 2413 931
rect 2430 914 2433 931
rect 2409 897 2433 914
rect 2409 880 2413 897
rect 2430 880 2433 897
rect 2409 863 2433 880
rect 2409 846 2413 863
rect 2430 846 2433 863
rect 2409 829 2433 846
rect 2409 812 2413 829
rect 2430 812 2433 829
rect 2409 795 2433 812
rect 2409 778 2413 795
rect 2430 778 2433 795
rect 2409 761 2433 778
rect 2409 744 2413 761
rect 2430 744 2433 761
rect 2409 727 2433 744
rect 2409 710 2413 727
rect 2430 710 2433 727
rect 2409 693 2433 710
rect 2409 676 2413 693
rect 2430 676 2433 693
rect 2409 659 2433 676
rect 2409 642 2413 659
rect 2430 642 2433 659
rect 2409 625 2433 642
rect 2409 608 2413 625
rect 2430 608 2433 625
rect 2409 591 2433 608
rect 2409 574 2413 591
rect 2430 574 2433 591
rect 2409 557 2433 574
rect 2409 540 2413 557
rect 2430 540 2433 557
rect 2409 523 2433 540
rect 2409 506 2413 523
rect 2430 506 2433 523
rect 2409 489 2433 506
rect 2409 472 2413 489
rect 2430 472 2433 489
rect 2409 455 2433 472
rect 2409 438 2413 455
rect 2430 438 2433 455
rect 2409 421 2433 438
rect 2409 404 2413 421
rect 2430 404 2433 421
rect 2409 387 2433 404
rect 2409 370 2413 387
rect 2430 370 2433 387
rect 2409 353 2433 370
rect 2409 336 2413 353
rect 2430 336 2433 353
rect 2409 319 2433 336
rect 2409 302 2413 319
rect 2430 302 2433 319
rect 2409 285 2433 302
rect 2409 268 2413 285
rect 2430 268 2433 285
rect 2409 251 2433 268
rect 2409 234 2413 251
rect 2430 234 2433 251
rect 2409 217 2433 234
rect 2409 200 2413 217
rect 2430 200 2433 217
rect 2409 183 2433 200
rect 2409 166 2413 183
rect 2430 166 2433 183
rect 2409 115 2433 166
rect 2455 1135 2479 1184
rect 2455 1118 2458 1135
rect 2475 1118 2479 1135
rect 2455 1101 2479 1118
rect 2455 1084 2458 1101
rect 2475 1084 2479 1101
rect 2455 1067 2479 1084
rect 2455 1050 2458 1067
rect 2475 1050 2479 1067
rect 2455 1033 2479 1050
rect 2455 1016 2458 1033
rect 2475 1016 2479 1033
rect 2455 999 2479 1016
rect 2455 982 2459 999
rect 2476 982 2479 999
rect 2455 965 2479 982
rect 2455 948 2459 965
rect 2476 948 2479 965
rect 2455 931 2479 948
rect 2455 914 2459 931
rect 2476 914 2479 931
rect 2455 897 2479 914
rect 2455 880 2459 897
rect 2476 880 2479 897
rect 2455 863 2479 880
rect 2455 846 2459 863
rect 2476 846 2479 863
rect 2455 829 2479 846
rect 2455 812 2459 829
rect 2476 812 2479 829
rect 2455 795 2479 812
rect 2455 778 2459 795
rect 2476 778 2479 795
rect 2455 761 2479 778
rect 2455 744 2459 761
rect 2476 744 2479 761
rect 2455 727 2479 744
rect 2455 710 2459 727
rect 2476 710 2479 727
rect 2455 693 2479 710
rect 2455 676 2459 693
rect 2476 676 2479 693
rect 2455 659 2479 676
rect 2455 642 2459 659
rect 2476 642 2479 659
rect 2455 625 2479 642
rect 2455 608 2459 625
rect 2476 608 2479 625
rect 2455 591 2479 608
rect 2455 574 2459 591
rect 2476 574 2479 591
rect 2455 557 2479 574
rect 2455 540 2459 557
rect 2476 540 2479 557
rect 2455 523 2479 540
rect 2455 506 2459 523
rect 2476 506 2479 523
rect 2455 489 2479 506
rect 2455 472 2459 489
rect 2476 472 2479 489
rect 2455 455 2479 472
rect 2455 438 2459 455
rect 2476 438 2479 455
rect 2455 421 2479 438
rect 2455 404 2459 421
rect 2476 404 2479 421
rect 2455 387 2479 404
rect 2455 370 2459 387
rect 2476 370 2479 387
rect 2455 353 2479 370
rect 2455 336 2459 353
rect 2476 336 2479 353
rect 2455 319 2479 336
rect 2455 302 2459 319
rect 2476 302 2479 319
rect 2455 285 2479 302
rect 2455 268 2459 285
rect 2476 268 2479 285
rect 2455 251 2479 268
rect 2455 234 2459 251
rect 2476 234 2479 251
rect 2455 217 2479 234
rect 2455 200 2459 217
rect 2476 200 2479 217
rect 2455 183 2479 200
rect 2455 166 2459 183
rect 2476 166 2479 183
rect 2455 158 2479 166
rect 2500 1137 2523 1145
rect 2500 1120 2503 1137
rect 2520 1120 2523 1137
rect 2500 1103 2523 1120
rect 2500 1086 2503 1103
rect 2520 1086 2523 1103
rect 2500 1069 2523 1086
rect 2500 1052 2503 1069
rect 2520 1052 2523 1069
rect 2500 1035 2523 1052
rect 2500 1018 2503 1035
rect 2520 1018 2523 1035
rect 2500 1001 2523 1018
rect 2500 984 2503 1001
rect 2520 984 2523 1001
rect 2500 967 2523 984
rect 2500 950 2503 967
rect 2520 950 2523 967
rect 2500 933 2523 950
rect 2500 916 2503 933
rect 2520 916 2523 933
rect 2500 899 2523 916
rect 2500 882 2503 899
rect 2520 882 2523 899
rect 2500 865 2523 882
rect 2500 848 2503 865
rect 2520 848 2523 865
rect 2500 831 2523 848
rect 2500 814 2503 831
rect 2520 814 2523 831
rect 2500 797 2523 814
rect 2500 780 2503 797
rect 2520 780 2523 797
rect 2500 763 2523 780
rect 2500 746 2503 763
rect 2520 746 2523 763
rect 2500 729 2523 746
rect 2500 712 2503 729
rect 2520 712 2523 729
rect 2500 695 2523 712
rect 2500 678 2503 695
rect 2520 678 2523 695
rect 2500 661 2523 678
rect 2500 644 2503 661
rect 2520 644 2523 661
rect 2500 627 2523 644
rect 2500 610 2503 627
rect 2520 610 2523 627
rect 2500 593 2523 610
rect 2500 576 2503 593
rect 2520 576 2523 593
rect 2500 559 2523 576
rect 2500 542 2503 559
rect 2520 542 2523 559
rect 2500 525 2523 542
rect 2500 508 2503 525
rect 2520 508 2523 525
rect 2500 491 2523 508
rect 2500 474 2503 491
rect 2520 474 2523 491
rect 2500 457 2523 474
rect 2500 440 2503 457
rect 2520 440 2523 457
rect 2500 423 2523 440
rect 2500 406 2503 423
rect 2520 406 2523 423
rect 2500 389 2523 406
rect 2500 372 2503 389
rect 2520 372 2523 389
rect 2500 355 2523 372
rect 2500 338 2503 355
rect 2520 338 2523 355
rect 2500 321 2523 338
rect 2500 304 2503 321
rect 2520 304 2523 321
rect 2500 287 2523 304
rect 2500 270 2503 287
rect 2520 270 2523 287
rect 2500 253 2523 270
rect 2500 236 2503 253
rect 2520 236 2523 253
rect 2500 219 2523 236
rect 2500 202 2503 219
rect 2520 202 2523 219
rect 2500 185 2523 202
rect 2500 168 2503 185
rect 2520 168 2523 185
rect 2500 115 2523 168
rect 2544 1135 2568 1184
rect 2544 1118 2547 1135
rect 2564 1118 2568 1135
rect 2544 1101 2568 1118
rect 2544 1084 2547 1101
rect 2564 1084 2568 1101
rect 2544 1067 2568 1084
rect 2544 1050 2547 1067
rect 2564 1050 2568 1067
rect 2544 1033 2568 1050
rect 2544 1016 2547 1033
rect 2564 1016 2568 1033
rect 2544 999 2568 1016
rect 2544 982 2548 999
rect 2565 982 2568 999
rect 2544 965 2568 982
rect 2544 948 2548 965
rect 2565 948 2568 965
rect 2544 931 2568 948
rect 2544 914 2548 931
rect 2565 914 2568 931
rect 2544 897 2568 914
rect 2544 880 2548 897
rect 2565 880 2568 897
rect 2544 863 2568 880
rect 2544 846 2548 863
rect 2565 846 2568 863
rect 2544 829 2568 846
rect 2544 812 2548 829
rect 2565 812 2568 829
rect 2544 795 2568 812
rect 2544 778 2548 795
rect 2565 778 2568 795
rect 2544 761 2568 778
rect 2544 744 2548 761
rect 2565 744 2568 761
rect 2544 727 2568 744
rect 2544 710 2548 727
rect 2565 710 2568 727
rect 2544 693 2568 710
rect 2544 676 2548 693
rect 2565 676 2568 693
rect 2544 659 2568 676
rect 2544 642 2548 659
rect 2565 642 2568 659
rect 2544 625 2568 642
rect 2544 608 2548 625
rect 2565 608 2568 625
rect 2544 591 2568 608
rect 2544 574 2548 591
rect 2565 574 2568 591
rect 2544 557 2568 574
rect 2544 540 2548 557
rect 2565 540 2568 557
rect 2544 523 2568 540
rect 2544 506 2548 523
rect 2565 506 2568 523
rect 2544 489 2568 506
rect 2544 472 2548 489
rect 2565 472 2568 489
rect 2544 455 2568 472
rect 2544 438 2548 455
rect 2565 438 2568 455
rect 2544 421 2568 438
rect 2544 404 2548 421
rect 2565 404 2568 421
rect 2544 387 2568 404
rect 2544 370 2548 387
rect 2565 370 2568 387
rect 2544 353 2568 370
rect 2544 336 2548 353
rect 2565 336 2568 353
rect 2544 319 2568 336
rect 2544 302 2548 319
rect 2565 302 2568 319
rect 2544 285 2568 302
rect 2544 268 2548 285
rect 2565 268 2568 285
rect 2544 251 2568 268
rect 2544 234 2548 251
rect 2565 234 2568 251
rect 2544 217 2568 234
rect 2544 200 2548 217
rect 2565 200 2568 217
rect 2544 183 2568 200
rect 2544 166 2548 183
rect 2565 166 2568 183
rect 2544 158 2568 166
rect 2589 1135 2613 1143
rect 2589 1118 2592 1135
rect 2609 1118 2613 1135
rect 2589 1101 2613 1118
rect 2589 1084 2592 1101
rect 2609 1084 2613 1101
rect 2589 1067 2613 1084
rect 2589 1050 2592 1067
rect 2609 1050 2613 1067
rect 2589 1033 2613 1050
rect 2589 1016 2592 1033
rect 2609 1016 2613 1033
rect 2589 999 2613 1016
rect 2589 982 2593 999
rect 2610 982 2613 999
rect 2589 965 2613 982
rect 2589 948 2593 965
rect 2610 948 2613 965
rect 2589 931 2613 948
rect 2589 914 2593 931
rect 2610 914 2613 931
rect 2589 897 2613 914
rect 2589 880 2593 897
rect 2610 880 2613 897
rect 2589 863 2613 880
rect 2589 846 2593 863
rect 2610 846 2613 863
rect 2589 829 2613 846
rect 2589 812 2593 829
rect 2610 812 2613 829
rect 2589 795 2613 812
rect 2589 778 2593 795
rect 2610 778 2613 795
rect 2589 761 2613 778
rect 2589 744 2593 761
rect 2610 744 2613 761
rect 2589 727 2613 744
rect 2589 710 2593 727
rect 2610 710 2613 727
rect 2589 693 2613 710
rect 2589 676 2593 693
rect 2610 676 2613 693
rect 2589 659 2613 676
rect 2589 642 2593 659
rect 2610 642 2613 659
rect 2589 625 2613 642
rect 2589 608 2593 625
rect 2610 608 2613 625
rect 2589 591 2613 608
rect 2589 574 2593 591
rect 2610 574 2613 591
rect 2589 557 2613 574
rect 2589 540 2593 557
rect 2610 540 2613 557
rect 2589 523 2613 540
rect 2589 506 2593 523
rect 2610 506 2613 523
rect 2589 489 2613 506
rect 2589 472 2593 489
rect 2610 472 2613 489
rect 2589 455 2613 472
rect 2589 438 2593 455
rect 2610 438 2613 455
rect 2589 421 2613 438
rect 2589 404 2593 421
rect 2610 404 2613 421
rect 2589 387 2613 404
rect 2589 370 2593 387
rect 2610 370 2613 387
rect 2589 353 2613 370
rect 2589 336 2593 353
rect 2610 336 2613 353
rect 2589 319 2613 336
rect 2589 302 2593 319
rect 2610 302 2613 319
rect 2589 285 2613 302
rect 2589 268 2593 285
rect 2610 268 2613 285
rect 2589 251 2613 268
rect 2589 234 2593 251
rect 2610 234 2613 251
rect 2589 217 2613 234
rect 2589 200 2593 217
rect 2610 200 2613 217
rect 2589 183 2613 200
rect 2589 166 2593 183
rect 2610 166 2613 183
rect 2589 115 2613 166
rect 2634 1135 2660 1184
rect 2634 1118 2637 1135
rect 2654 1118 2660 1135
rect 2634 1101 2660 1118
rect 2634 1084 2637 1101
rect 2654 1084 2660 1101
rect 2634 1067 2660 1084
rect 2634 1050 2637 1067
rect 2654 1050 2660 1067
rect 2634 1033 2660 1050
rect 2634 1016 2637 1033
rect 2654 1016 2660 1033
rect 2634 999 2660 1016
rect 2634 982 2638 999
rect 2655 982 2660 999
rect 2634 965 2660 982
rect 2634 948 2638 965
rect 2655 948 2660 965
rect 2634 931 2660 948
rect 2634 914 2638 931
rect 2655 914 2660 931
rect 2634 897 2660 914
rect 2634 880 2638 897
rect 2655 880 2660 897
rect 2634 863 2660 880
rect 2634 846 2638 863
rect 2655 846 2660 863
rect 2634 829 2660 846
rect 2634 812 2638 829
rect 2655 812 2660 829
rect 2634 795 2660 812
rect 2634 778 2638 795
rect 2655 778 2660 795
rect 2634 761 2660 778
rect 2634 744 2638 761
rect 2655 744 2660 761
rect 2634 727 2660 744
rect 2634 710 2638 727
rect 2655 710 2660 727
rect 2634 693 2660 710
rect 2634 676 2638 693
rect 2655 676 2660 693
rect 2634 659 2660 676
rect 2634 642 2638 659
rect 2655 642 2660 659
rect 2634 625 2660 642
rect 2634 608 2638 625
rect 2655 608 2660 625
rect 2634 591 2660 608
rect 2634 574 2638 591
rect 2655 574 2660 591
rect 2634 557 2660 574
rect 2634 540 2638 557
rect 2655 540 2660 557
rect 2634 523 2660 540
rect 2634 506 2638 523
rect 2655 506 2660 523
rect 2634 489 2660 506
rect 2634 472 2638 489
rect 2655 472 2660 489
rect 2634 455 2660 472
rect 2634 438 2638 455
rect 2655 438 2660 455
rect 2634 421 2660 438
rect 2634 404 2638 421
rect 2655 404 2660 421
rect 2634 387 2660 404
rect 2634 370 2638 387
rect 2655 370 2660 387
rect 2634 353 2660 370
rect 2634 336 2638 353
rect 2655 336 2660 353
rect 2634 319 2660 336
rect 2634 302 2638 319
rect 2655 302 2660 319
rect 2634 285 2660 302
rect 2634 268 2638 285
rect 2655 268 2660 285
rect 2634 251 2660 268
rect 2634 234 2638 251
rect 2655 234 2660 251
rect 2634 217 2660 234
rect 2634 200 2638 217
rect 2655 200 2660 217
rect 2634 183 2660 200
rect 2634 166 2638 183
rect 2655 166 2660 183
rect 2634 158 2660 166
rect -17 112 2613 115
rect -17 111 983 112
rect -17 110 641 111
rect -17 93 -9 110
rect 8 109 196 110
rect 8 93 25 109
rect -17 92 25 93
rect 42 92 59 109
rect 76 108 128 109
rect 76 92 94 108
rect -17 91 94 92
rect 111 92 128 108
rect 145 92 162 109
rect 179 93 196 109
rect 213 93 230 110
rect 247 93 265 110
rect 282 93 299 110
rect 316 109 470 110
rect 316 108 367 109
rect 316 93 333 108
rect 179 92 333 93
rect 111 91 333 92
rect 350 92 367 108
rect 384 92 401 109
rect 418 92 436 109
rect 453 93 470 109
rect 487 93 504 110
rect 521 93 538 110
rect 555 93 572 110
rect 589 93 607 110
rect 624 94 641 110
rect 658 110 812 111
rect 658 94 675 110
rect 624 93 675 94
rect 692 93 709 110
rect 726 93 743 110
rect 760 93 778 110
rect 795 94 812 110
rect 829 94 846 111
rect 863 94 880 111
rect 897 94 914 111
rect 931 94 949 111
rect 966 95 983 111
rect 1000 111 1256 112
rect 1000 95 1017 111
rect 966 94 1017 95
rect 1034 94 1051 111
rect 1068 94 1085 111
rect 1102 94 1120 111
rect 1137 94 1154 111
rect 1171 94 1188 111
rect 1205 94 1222 111
rect 1239 95 1256 111
rect 1273 111 1325 112
rect 1273 95 1291 111
rect 1239 94 1291 95
rect 1308 95 1325 111
rect 1342 110 1393 112
rect 1342 95 1359 110
rect 1308 94 1359 95
rect 795 93 1359 94
rect 1376 95 1393 110
rect 1410 111 1804 112
rect 1410 95 1427 111
rect 1376 94 1427 95
rect 1444 94 1462 111
rect 1479 94 1496 111
rect 1513 110 1633 111
rect 1513 94 1530 110
rect 1376 93 1530 94
rect 1547 93 1564 110
rect 1581 93 1599 110
rect 1616 94 1633 110
rect 1650 94 1667 111
rect 1684 94 1701 111
rect 1718 94 1735 111
rect 1752 94 1770 111
rect 1787 95 1804 111
rect 1821 111 1872 112
rect 1821 95 1838 111
rect 1787 94 1838 95
rect 1855 95 1872 111
rect 1889 111 1941 112
rect 1889 95 1906 111
rect 1855 94 1906 95
rect 1923 95 1941 111
rect 1958 111 2284 112
rect 1958 95 1976 111
rect 1923 94 1976 95
rect 1993 110 2079 111
rect 1993 94 2010 110
rect 1616 93 2010 94
rect 2027 93 2044 110
rect 2061 94 2079 110
rect 2096 94 2113 111
rect 2130 94 2147 111
rect 2164 94 2181 111
rect 2198 94 2215 111
rect 2232 94 2250 111
rect 2267 95 2284 111
rect 2301 111 2352 112
rect 2301 95 2318 111
rect 2267 94 2318 95
rect 2335 95 2352 111
rect 2369 111 2421 112
rect 2369 95 2386 111
rect 2335 94 2386 95
rect 2403 95 2421 111
rect 2438 111 2613 112
rect 2438 95 2455 111
rect 2403 94 2455 95
rect 2472 94 2489 111
rect 2506 110 2613 111
rect 2506 94 2523 110
rect 2061 93 2523 94
rect 2540 93 2558 110
rect 2575 108 2613 110
rect 2575 93 2592 108
rect 453 92 2592 93
rect 350 91 2592 92
rect 2609 91 2613 108
rect -17 83 2613 91
<< viali >>
rect -79 1203 -62 1220
rect -43 1203 -26 1220
rect -7 1202 10 1219
rect 29 1202 46 1219
rect 65 1202 82 1219
rect 101 1202 118 1219
rect 137 1202 154 1219
rect 173 1202 190 1219
rect 209 1201 226 1218
rect 245 1201 262 1218
rect 281 1201 298 1218
rect 317 1201 334 1218
rect 354 1201 371 1218
rect 390 1201 407 1218
rect 426 1200 443 1217
rect 462 1200 479 1217
rect 498 1200 515 1217
rect 534 1200 551 1217
rect 570 1200 587 1217
rect 606 1200 623 1217
rect 642 1199 659 1216
rect 678 1199 695 1216
rect 714 1199 731 1216
rect 750 1199 767 1216
rect 787 1201 804 1218
rect 823 1201 840 1218
rect 859 1201 876 1218
rect 896 1201 913 1218
rect 932 1201 949 1218
rect 968 1200 985 1217
rect 1004 1200 1021 1217
rect 1040 1200 1057 1217
rect 1076 1200 1093 1217
rect 1112 1200 1129 1217
rect 1148 1200 1165 1217
rect 1185 1202 1202 1219
rect 1221 1202 1238 1219
rect 1257 1202 1274 1219
rect 1294 1202 1311 1219
rect 1330 1202 1347 1219
rect 1366 1201 1383 1218
rect 1402 1201 1419 1218
rect 1438 1201 1455 1218
rect 1474 1201 1491 1218
rect 1510 1201 1527 1218
rect 1546 1201 1563 1218
rect 1582 1202 1599 1219
rect 1618 1202 1635 1219
rect 1654 1202 1671 1219
rect 1691 1202 1708 1219
rect 1727 1202 1744 1219
rect 1763 1201 1780 1218
rect 1799 1201 1816 1218
rect 1835 1201 1852 1218
rect 1871 1201 1888 1218
rect 1907 1201 1924 1218
rect 1943 1201 1960 1218
rect 1979 1202 1996 1219
rect 2015 1202 2032 1219
rect 2051 1202 2068 1219
rect 2088 1202 2105 1219
rect 2124 1202 2141 1219
rect 2160 1201 2177 1218
rect 2196 1201 2213 1218
rect 2232 1201 2249 1218
rect 2268 1201 2285 1218
rect 2304 1201 2321 1218
rect 2340 1201 2357 1218
rect 2376 1202 2393 1219
rect 2412 1202 2429 1219
rect 2448 1201 2465 1218
rect 2484 1201 2501 1218
rect 2525 1201 2542 1218
rect 2561 1201 2578 1218
rect 2601 1201 2618 1218
rect 2642 1201 2659 1218
rect -9 93 8 110
rect 59 92 76 109
rect 128 92 145 109
rect 196 93 213 110
rect 265 93 282 110
rect 333 91 350 108
rect 401 92 418 109
rect 470 93 487 110
rect 538 93 555 110
rect 607 93 624 110
rect 675 93 692 110
rect 743 93 760 110
rect 812 94 829 111
rect 880 94 897 111
rect 949 94 966 111
rect 1017 94 1034 111
rect 1085 94 1102 111
rect 1154 94 1171 111
rect 1222 94 1239 111
rect 1291 94 1308 111
rect 1359 93 1376 110
rect 1427 94 1444 111
rect 1496 94 1513 111
rect 1564 93 1581 110
rect 1633 94 1650 111
rect 1701 94 1718 111
rect 1770 94 1787 111
rect 1838 94 1855 111
rect 1906 94 1923 111
rect 1976 94 1993 111
rect 2044 93 2061 110
rect 2113 94 2130 111
rect 2181 94 2198 111
rect 2250 94 2267 111
rect 2318 94 2335 111
rect 2386 94 2403 111
rect 2455 94 2472 111
rect 2523 93 2540 110
rect 2592 91 2609 108
<< metal1 >>
rect -85 1220 2677 1253
rect -85 1203 -79 1220
rect -62 1203 -43 1220
rect -26 1219 2677 1220
rect -26 1203 -7 1219
rect -85 1202 -7 1203
rect 10 1202 29 1219
rect 46 1202 65 1219
rect 82 1202 101 1219
rect 118 1202 137 1219
rect 154 1202 173 1219
rect 190 1218 1185 1219
rect 190 1202 209 1218
rect -85 1201 209 1202
rect 226 1201 245 1218
rect 262 1201 281 1218
rect 298 1201 317 1218
rect 334 1201 354 1218
rect 371 1201 390 1218
rect 407 1217 787 1218
rect 407 1201 426 1217
rect -85 1200 426 1201
rect 443 1200 462 1217
rect 479 1200 498 1217
rect 515 1200 534 1217
rect 551 1200 570 1217
rect 587 1200 606 1217
rect 623 1216 787 1217
rect 623 1200 642 1216
rect -85 1199 642 1200
rect 659 1199 678 1216
rect 695 1199 714 1216
rect 731 1199 750 1216
rect 767 1201 787 1216
rect 804 1201 823 1218
rect 840 1201 859 1218
rect 876 1201 896 1218
rect 913 1201 932 1218
rect 949 1217 1185 1218
rect 949 1201 968 1217
rect 767 1200 968 1201
rect 985 1200 1004 1217
rect 1021 1200 1040 1217
rect 1057 1200 1076 1217
rect 1093 1200 1112 1217
rect 1129 1200 1148 1217
rect 1165 1202 1185 1217
rect 1202 1202 1221 1219
rect 1238 1202 1257 1219
rect 1274 1202 1294 1219
rect 1311 1202 1330 1219
rect 1347 1218 1582 1219
rect 1347 1202 1366 1218
rect 1165 1201 1366 1202
rect 1383 1201 1402 1218
rect 1419 1201 1438 1218
rect 1455 1201 1474 1218
rect 1491 1201 1510 1218
rect 1527 1201 1546 1218
rect 1563 1202 1582 1218
rect 1599 1202 1618 1219
rect 1635 1202 1654 1219
rect 1671 1202 1691 1219
rect 1708 1202 1727 1219
rect 1744 1218 1979 1219
rect 1744 1202 1763 1218
rect 1563 1201 1763 1202
rect 1780 1201 1799 1218
rect 1816 1201 1835 1218
rect 1852 1201 1871 1218
rect 1888 1201 1907 1218
rect 1924 1201 1943 1218
rect 1960 1202 1979 1218
rect 1996 1202 2015 1219
rect 2032 1202 2051 1219
rect 2068 1202 2088 1219
rect 2105 1202 2124 1219
rect 2141 1218 2376 1219
rect 2141 1202 2160 1218
rect 1960 1201 2160 1202
rect 2177 1201 2196 1218
rect 2213 1201 2232 1218
rect 2249 1201 2268 1218
rect 2285 1201 2304 1218
rect 2321 1201 2340 1218
rect 2357 1202 2376 1218
rect 2393 1202 2412 1219
rect 2429 1218 2677 1219
rect 2429 1202 2448 1218
rect 2357 1201 2448 1202
rect 2465 1201 2484 1218
rect 2501 1201 2525 1218
rect 2542 1201 2561 1218
rect 2578 1201 2601 1218
rect 2618 1201 2642 1218
rect 2659 1201 2677 1218
rect 1165 1200 2677 1201
rect 767 1199 2677 1200
rect -85 1195 2677 1199
rect -85 1194 2660 1195
rect -17 111 2613 114
rect -17 110 812 111
rect -17 93 -9 110
rect 8 109 196 110
rect 8 93 59 109
rect -17 92 59 93
rect 76 92 128 109
rect 145 93 196 109
rect 213 93 265 110
rect 282 109 470 110
rect 282 108 401 109
rect 282 93 333 108
rect 145 92 333 93
rect -17 91 333 92
rect 350 92 401 108
rect 418 93 470 109
rect 487 93 538 110
rect 555 93 607 110
rect 624 93 675 110
rect 692 93 743 110
rect 760 94 812 110
rect 829 94 880 111
rect 897 94 949 111
rect 966 94 1017 111
rect 1034 94 1085 111
rect 1102 94 1154 111
rect 1171 94 1222 111
rect 1239 94 1291 111
rect 1308 110 1427 111
rect 1308 94 1359 110
rect 760 93 1359 94
rect 1376 94 1427 110
rect 1444 94 1496 111
rect 1513 110 1633 111
rect 1513 94 1564 110
rect 1376 93 1564 94
rect 1581 94 1633 110
rect 1650 94 1701 111
rect 1718 94 1770 111
rect 1787 94 1838 111
rect 1855 94 1906 111
rect 1923 94 1976 111
rect 1993 110 2113 111
rect 1993 94 2044 110
rect 1581 93 2044 94
rect 2061 94 2113 110
rect 2130 94 2181 111
rect 2198 94 2250 111
rect 2267 94 2318 111
rect 2335 94 2386 111
rect 2403 94 2455 111
rect 2472 110 2613 111
rect 2472 94 2523 110
rect 2061 93 2523 94
rect 2540 108 2613 110
rect 2540 93 2592 108
rect 418 92 2592 93
rect 350 91 2592 92
rect 2609 91 2613 108
rect -17 62 2613 91
<< labels >>
rlabel metal1 -85 1253 2677 1253 1 VP
rlabel metal1 -17 62 2613 62 5 VN
<< end >>
